library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"fcf2c487",
    12 => x"86c0c64e",
    13 => x"49fcf2c4",
    14 => x"48e4f9c3",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087f4eb",
    19 => x"1e87fc98",
    20 => x"48121e72",
    21 => x"87c40211",
    22 => x"87f60288",
    23 => x"4f264a26",
    24 => x"731e721e",
    25 => x"1148121e",
    26 => x"4b87ca02",
    27 => x"9b98dfc3",
    28 => x"f0028873",
    29 => x"264b2687",
    30 => x"1e4f264a",
    31 => x"1e721e73",
    32 => x"ca048bc1",
    33 => x"11481287",
    34 => x"8887c402",
    35 => x"2687f102",
    36 => x"264b264a",
    37 => x"1e741e4f",
    38 => x"1e721e73",
    39 => x"d0048bc1",
    40 => x"11481287",
    41 => x"4c87ca02",
    42 => x"9c98dfc3",
    43 => x"eb028874",
    44 => x"264a2687",
    45 => x"264c264b",
    46 => x"48731e4f",
    47 => x"02a97381",
    48 => x"531287c5",
    49 => x"2687f605",
    50 => x"66c41e4f",
    51 => x"1248714a",
    52 => x"87fb0551",
    53 => x"731e4f26",
    54 => x"a9738148",
    55 => x"f9537205",
    56 => x"0e4f2687",
    57 => x"5d5c5b5e",
    58 => x"7186f40e",
    59 => x"48a6c44d",
    60 => x"66dc78c0",
    61 => x"48a6c84b",
    62 => x"971578c0",
    63 => x"026e977e",
    64 => x"1387f0c0",
    65 => x"da029c4c",
    66 => x"4a6e9787",
    67 => x"aab74974",
    68 => x"c887c905",
    69 => x"78c148a6",
    70 => x"87c24cc0",
    71 => x"9c744c13",
    72 => x"c887e605",
    73 => x"87cb0266",
    74 => x"c14866c4",
    75 => x"58a6c880",
    76 => x"c487fffe",
    77 => x"8ef44866",
    78 => x"4c264d26",
    79 => x"4f264b26",
    80 => x"c14a711e",
    81 => x"04aab7c1",
    82 => x"c6c187d9",
    83 => x"d201aab7",
    84 => x"4866c487",
    85 => x"ca05a8d0",
    86 => x"c0497287",
    87 => x"487189f7",
    88 => x"c187ecc0",
    89 => x"04aab7e1",
    90 => x"e6c187d8",
    91 => x"d101aab7",
    92 => x"4866c487",
    93 => x"c905a8d0",
    94 => x"c1497287",
    95 => x"487189d7",
    96 => x"f0c087cd",
    97 => x"aab7c98a",
    98 => x"ff87c206",
    99 => x"2648724a",
   100 => x"5b5e0e4f",
   101 => x"f80e5d5c",
   102 => x"c47e7186",
   103 => x"78c048a6",
   104 => x"a7f9c14c",
   105 => x"4966c41e",
   106 => x"c487f8fc",
   107 => x"6e497086",
   108 => x"9783714b",
   109 => x"edc0496b",
   110 => x"87c605a9",
   111 => x"c148a6c4",
   112 => x"66d88378",
   113 => x"d887c502",
   114 => x"0b7b0b66",
   115 => x"d3056b97",
   116 => x"0266c487",
   117 => x"4a7487c7",
   118 => x"c28a0ac0",
   119 => x"724a7487",
   120 => x"87efc048",
   121 => x"131e66dc",
   122 => x"87d4fd49",
   123 => x"4d7086c4",
   124 => x"03adb7c0",
   125 => x"66c487d4",
   126 => x"7487c902",
   127 => x"8808c048",
   128 => x"87c27e70",
   129 => x"486e7e74",
   130 => x"66dc87c9",
   131 => x"4ca47594",
   132 => x"f887effe",
   133 => x"264d268e",
   134 => x"264b264c",
   135 => x"1e00204f",
   136 => x"9a721e73",
   137 => x"87e7c002",
   138 => x"4bc148c0",
   139 => x"d106a972",
   140 => x"06827287",
   141 => x"837387c9",
   142 => x"f401a972",
   143 => x"c187c387",
   144 => x"a9723ab2",
   145 => x"80738903",
   146 => x"2b2ac107",
   147 => x"2687f305",
   148 => x"1e4f264b",
   149 => x"4dc41e75",
   150 => x"04a1b771",
   151 => x"81c1b9ff",
   152 => x"7207bdc3",
   153 => x"ff04a2b7",
   154 => x"c182c1ba",
   155 => x"eefe07bd",
   156 => x"042dc187",
   157 => x"80c1b8ff",
   158 => x"ff042d07",
   159 => x"0781c1b9",
   160 => x"4f264d26",
   161 => x"ff48111e",
   162 => x"c47808d4",
   163 => x"88c14866",
   164 => x"7058a6c8",
   165 => x"87ed0598",
   166 => x"ff1e4f26",
   167 => x"ffc348d4",
   168 => x"c4516878",
   169 => x"88c14866",
   170 => x"7058a6c8",
   171 => x"87eb0598",
   172 => x"731e4f26",
   173 => x"4bd4ff1e",
   174 => x"6b7bffc3",
   175 => x"7bffc34a",
   176 => x"32c8496b",
   177 => x"ffc3b172",
   178 => x"c84a6b7b",
   179 => x"c3b27131",
   180 => x"496b7bff",
   181 => x"b17232c8",
   182 => x"87c44871",
   183 => x"4c264d26",
   184 => x"4f264b26",
   185 => x"5c5b5e0e",
   186 => x"4a710e5d",
   187 => x"724cd4ff",
   188 => x"99ffc349",
   189 => x"f9c37c71",
   190 => x"c805bfe4",
   191 => x"4866d087",
   192 => x"a6d430c9",
   193 => x"4966d058",
   194 => x"ffc329d8",
   195 => x"d07c7199",
   196 => x"29d04966",
   197 => x"7199ffc3",
   198 => x"4966d07c",
   199 => x"ffc329c8",
   200 => x"d07c7199",
   201 => x"ffc34966",
   202 => x"727c7199",
   203 => x"c329d049",
   204 => x"7c7199ff",
   205 => x"f0c94b6c",
   206 => x"ffc34dff",
   207 => x"87d005ab",
   208 => x"6c7cffc3",
   209 => x"028dc14b",
   210 => x"ffc387c6",
   211 => x"87f002ab",
   212 => x"c7fe4873",
   213 => x"49c01e87",
   214 => x"c348d4ff",
   215 => x"81c178ff",
   216 => x"a9b7c8c3",
   217 => x"2687f104",
   218 => x"1e731e4f",
   219 => x"f8c487e7",
   220 => x"1ec04bdf",
   221 => x"c1f0ffc0",
   222 => x"e7fd49f7",
   223 => x"c186c487",
   224 => x"eac005a8",
   225 => x"48d4ff87",
   226 => x"c178ffc3",
   227 => x"c0c0c0c0",
   228 => x"e1c01ec0",
   229 => x"49e9c1f0",
   230 => x"c487c9fd",
   231 => x"05987086",
   232 => x"d4ff87ca",
   233 => x"78ffc348",
   234 => x"87cb48c1",
   235 => x"c187e6fe",
   236 => x"fdfe058b",
   237 => x"fc48c087",
   238 => x"731e87e6",
   239 => x"48d4ff1e",
   240 => x"d378ffc3",
   241 => x"c01ec04b",
   242 => x"c1c1f0ff",
   243 => x"87d4fc49",
   244 => x"987086c4",
   245 => x"ff87ca05",
   246 => x"ffc348d4",
   247 => x"cb48c178",
   248 => x"87f1fd87",
   249 => x"ff058bc1",
   250 => x"48c087db",
   251 => x"0e87f1fb",
   252 => x"0e5c5b5e",
   253 => x"fd4cd4ff",
   254 => x"eac687db",
   255 => x"f0e1c01e",
   256 => x"fb49c8c1",
   257 => x"86c487de",
   258 => x"c802a8c1",
   259 => x"87eafe87",
   260 => x"e2c148c0",
   261 => x"87dafa87",
   262 => x"ffcf4970",
   263 => x"eac699ff",
   264 => x"87c802a9",
   265 => x"c087d3fe",
   266 => x"87cbc148",
   267 => x"c07cffc3",
   268 => x"f4fc4bf1",
   269 => x"02987087",
   270 => x"c087ebc0",
   271 => x"f0ffc01e",
   272 => x"fa49fac1",
   273 => x"86c487de",
   274 => x"d9059870",
   275 => x"7cffc387",
   276 => x"ffc3496c",
   277 => x"7c7c7c7c",
   278 => x"0299c0c1",
   279 => x"48c187c4",
   280 => x"48c087d5",
   281 => x"abc287d1",
   282 => x"c087c405",
   283 => x"c187c848",
   284 => x"fdfe058b",
   285 => x"f948c087",
   286 => x"731e87e4",
   287 => x"e4f9c31e",
   288 => x"c778c148",
   289 => x"48d0ff4b",
   290 => x"c8fb78c2",
   291 => x"48d0ff87",
   292 => x"1ec078c3",
   293 => x"c1d0e5c0",
   294 => x"c7f949c0",
   295 => x"c186c487",
   296 => x"87c105a8",
   297 => x"05abc24b",
   298 => x"48c087c5",
   299 => x"c187f9c0",
   300 => x"d0ff058b",
   301 => x"87f7fc87",
   302 => x"58e8f9c3",
   303 => x"cd059870",
   304 => x"c01ec187",
   305 => x"d0c1f0ff",
   306 => x"87d8f849",
   307 => x"d4ff86c4",
   308 => x"78ffc348",
   309 => x"c387e0c4",
   310 => x"ff58ecf9",
   311 => x"78c248d0",
   312 => x"c348d4ff",
   313 => x"48c178ff",
   314 => x"0e87f5f7",
   315 => x"5d5c5b5e",
   316 => x"c34a710e",
   317 => x"d4ff4dff",
   318 => x"ff7c754c",
   319 => x"c3c448d0",
   320 => x"727c7578",
   321 => x"f0ffc01e",
   322 => x"f749d8c1",
   323 => x"86c487d6",
   324 => x"c5029870",
   325 => x"c048c087",
   326 => x"7c7587f0",
   327 => x"c87cfec3",
   328 => x"66d41ec0",
   329 => x"87dcf549",
   330 => x"7c7586c4",
   331 => x"7c757c75",
   332 => x"4be0dad8",
   333 => x"496c7c75",
   334 => x"87c50599",
   335 => x"f3058bc1",
   336 => x"ff7c7587",
   337 => x"78c248d0",
   338 => x"cff648c1",
   339 => x"d4ff1e87",
   340 => x"48d0ff4a",
   341 => x"c378d1c4",
   342 => x"89c17aff",
   343 => x"2687f805",
   344 => x"1e731e4f",
   345 => x"eec54b71",
   346 => x"ff4adfcd",
   347 => x"ffc348d4",
   348 => x"c3486878",
   349 => x"c502a8fe",
   350 => x"058ac187",
   351 => x"9a7287ed",
   352 => x"c087c505",
   353 => x"87eac048",
   354 => x"cc029b73",
   355 => x"1e66c887",
   356 => x"c5f44973",
   357 => x"c686c487",
   358 => x"4966c887",
   359 => x"ff87eefe",
   360 => x"ffc348d4",
   361 => x"9b737878",
   362 => x"ff87c505",
   363 => x"78d048d0",
   364 => x"ebf448c1",
   365 => x"1e731e87",
   366 => x"4bc04a71",
   367 => x"c348d4ff",
   368 => x"d0ff78ff",
   369 => x"78c3c448",
   370 => x"c348d4ff",
   371 => x"1e7278ff",
   372 => x"c1f0ffc0",
   373 => x"cbf449d1",
   374 => x"7086c487",
   375 => x"87cd0598",
   376 => x"cc1ec0c8",
   377 => x"f8fd4966",
   378 => x"7086c487",
   379 => x"48d0ff4b",
   380 => x"487378c2",
   381 => x"0e87e9f3",
   382 => x"5d5c5b5e",
   383 => x"c01ec00e",
   384 => x"c9c1f0ff",
   385 => x"87dcf349",
   386 => x"f9c31ed2",
   387 => x"d0fd49ec",
   388 => x"c086c887",
   389 => x"d284c14c",
   390 => x"f804acb7",
   391 => x"ecf9c387",
   392 => x"c349bf97",
   393 => x"c0c199c0",
   394 => x"e7c005a9",
   395 => x"f3f9c387",
   396 => x"d049bf97",
   397 => x"f4f9c331",
   398 => x"c84abf97",
   399 => x"c3b17232",
   400 => x"bf97f5f9",
   401 => x"4c71b14a",
   402 => x"ffffffcf",
   403 => x"ca84c19c",
   404 => x"87e7c134",
   405 => x"97f5f9c3",
   406 => x"31c149bf",
   407 => x"f9c399c6",
   408 => x"4abf97f6",
   409 => x"722ab7c7",
   410 => x"f1f9c3b1",
   411 => x"4d4abf97",
   412 => x"f9c39dcf",
   413 => x"4abf97f2",
   414 => x"32ca9ac3",
   415 => x"97f3f9c3",
   416 => x"33c24bbf",
   417 => x"f9c3b273",
   418 => x"4bbf97f4",
   419 => x"c69bc0c3",
   420 => x"b2732bb7",
   421 => x"48c181c2",
   422 => x"49703071",
   423 => x"307548c1",
   424 => x"4c724d70",
   425 => x"947184c1",
   426 => x"adb7c0c8",
   427 => x"c187cc06",
   428 => x"c82db734",
   429 => x"01adb7c0",
   430 => x"7487f4ff",
   431 => x"87dcf048",
   432 => x"5c5b5e0e",
   433 => x"86f80e5d",
   434 => x"48d2c2c4",
   435 => x"fac378c0",
   436 => x"49c01eca",
   437 => x"c487defb",
   438 => x"05987086",
   439 => x"48c087c5",
   440 => x"c087cec9",
   441 => x"c07ec14d",
   442 => x"49bff9fe",
   443 => x"4ac0fbc3",
   444 => x"e64bc871",
   445 => x"987087c5",
   446 => x"c087c205",
   447 => x"f5fec07e",
   448 => x"fbc349bf",
   449 => x"c8714adc",
   450 => x"87efe54b",
   451 => x"c2059870",
   452 => x"6e7ec087",
   453 => x"87fdc002",
   454 => x"bfd0c1c4",
   455 => x"c8c2c44d",
   456 => x"487ebf9f",
   457 => x"a8ead6c5",
   458 => x"c487c705",
   459 => x"4dbfd0c1",
   460 => x"486e87ce",
   461 => x"a8d5e9ca",
   462 => x"c087c502",
   463 => x"87f1c748",
   464 => x"1ecafac3",
   465 => x"ecf94975",
   466 => x"7086c487",
   467 => x"87c50598",
   468 => x"dcc748c0",
   469 => x"f5fec087",
   470 => x"fbc349bf",
   471 => x"c8714adc",
   472 => x"87d7e44b",
   473 => x"c8059870",
   474 => x"d2c2c487",
   475 => x"da78c148",
   476 => x"f9fec087",
   477 => x"fbc349bf",
   478 => x"c8714ac0",
   479 => x"87fbe34b",
   480 => x"c0029870",
   481 => x"48c087c5",
   482 => x"c487e6c6",
   483 => x"bf97c8c2",
   484 => x"a9d5c149",
   485 => x"87cdc005",
   486 => x"97c9c2c4",
   487 => x"eac249bf",
   488 => x"c5c002a9",
   489 => x"c648c087",
   490 => x"fac387c7",
   491 => x"7ebf97ca",
   492 => x"a8e9c348",
   493 => x"87cec002",
   494 => x"ebc3486e",
   495 => x"c5c002a8",
   496 => x"c548c087",
   497 => x"fac387eb",
   498 => x"49bf97d5",
   499 => x"ccc00599",
   500 => x"d6fac387",
   501 => x"c249bf97",
   502 => x"c5c002a9",
   503 => x"c548c087",
   504 => x"fac387cf",
   505 => x"48bf97d7",
   506 => x"58cec2c4",
   507 => x"c1484c70",
   508 => x"d2c2c488",
   509 => x"d8fac358",
   510 => x"7549bf97",
   511 => x"d9fac381",
   512 => x"c84abf97",
   513 => x"7ea17232",
   514 => x"48dfc6c4",
   515 => x"fac3786e",
   516 => x"48bf97da",
   517 => x"c458a6c8",
   518 => x"02bfd2c2",
   519 => x"c087d4c2",
   520 => x"49bff5fe",
   521 => x"4adcfbc3",
   522 => x"e14bc871",
   523 => x"987087cd",
   524 => x"87c5c002",
   525 => x"f8c348c0",
   526 => x"cac2c487",
   527 => x"c6c44cbf",
   528 => x"fac35cf3",
   529 => x"49bf97ef",
   530 => x"fac331c8",
   531 => x"4abf97ee",
   532 => x"fac349a1",
   533 => x"4abf97f0",
   534 => x"a17232d0",
   535 => x"f1fac349",
   536 => x"d84abf97",
   537 => x"49a17232",
   538 => x"c49166c4",
   539 => x"81bfdfc6",
   540 => x"59e7c6c4",
   541 => x"97f7fac3",
   542 => x"32c84abf",
   543 => x"97f6fac3",
   544 => x"4aa24bbf",
   545 => x"97f8fac3",
   546 => x"33d04bbf",
   547 => x"c34aa273",
   548 => x"bf97f9fa",
   549 => x"d89bcf4b",
   550 => x"4aa27333",
   551 => x"5aebc6c4",
   552 => x"bfe7c6c4",
   553 => x"748ac24a",
   554 => x"ebc6c492",
   555 => x"78a17248",
   556 => x"c387cac1",
   557 => x"bf97dcfa",
   558 => x"c331c849",
   559 => x"bf97dbfa",
   560 => x"c449a14a",
   561 => x"c459dac2",
   562 => x"49bfd6c2",
   563 => x"ffc731c5",
   564 => x"c429c981",
   565 => x"c359f3c6",
   566 => x"bf97e1fa",
   567 => x"c332c84a",
   568 => x"bf97e0fa",
   569 => x"c44aa24b",
   570 => x"826e9266",
   571 => x"5aefc6c4",
   572 => x"48e7c6c4",
   573 => x"c6c478c0",
   574 => x"a17248e3",
   575 => x"f3c6c478",
   576 => x"e7c6c448",
   577 => x"c6c478bf",
   578 => x"c6c448f7",
   579 => x"c478bfeb",
   580 => x"02bfd2c2",
   581 => x"7487c9c0",
   582 => x"7030c448",
   583 => x"87c9c07e",
   584 => x"bfefc6c4",
   585 => x"7030c448",
   586 => x"d6c2c47e",
   587 => x"c1786e48",
   588 => x"268ef848",
   589 => x"264c264d",
   590 => x"0e4f264b",
   591 => x"5d5c5b5e",
   592 => x"c44a710e",
   593 => x"02bfd2c2",
   594 => x"4b7287cb",
   595 => x"4c722bc7",
   596 => x"c99cffc1",
   597 => x"c84b7287",
   598 => x"c34c722b",
   599 => x"c6c49cff",
   600 => x"c083bfdf",
   601 => x"abbff1fe",
   602 => x"c087d902",
   603 => x"c35bf5fe",
   604 => x"731ecafa",
   605 => x"87fdf049",
   606 => x"987086c4",
   607 => x"c087c505",
   608 => x"87e6c048",
   609 => x"bfd2c2c4",
   610 => x"7487d202",
   611 => x"c391c449",
   612 => x"6981cafa",
   613 => x"ffffcf4d",
   614 => x"cb9dffff",
   615 => x"c2497487",
   616 => x"cafac391",
   617 => x"4d699f81",
   618 => x"c6fe4875",
   619 => x"5b5e0e87",
   620 => x"1e0e5d5c",
   621 => x"1ec04d71",
   622 => x"dcd049c1",
   623 => x"7086c487",
   624 => x"c1029c4c",
   625 => x"c2c487c2",
   626 => x"49754ada",
   627 => x"87d0daff",
   628 => x"c0029870",
   629 => x"4a7487f2",
   630 => x"4bcb4975",
   631 => x"87f5daff",
   632 => x"c0029870",
   633 => x"1ec087e2",
   634 => x"c7029c74",
   635 => x"48a6c487",
   636 => x"87c578c0",
   637 => x"c148a6c4",
   638 => x"4966c478",
   639 => x"c487dacf",
   640 => x"9c4c7086",
   641 => x"87fefe05",
   642 => x"fc264874",
   643 => x"5e0e87e5",
   644 => x"0e5d5c5b",
   645 => x"9b4b711e",
   646 => x"c087c505",
   647 => x"87e5c148",
   648 => x"c04da3c8",
   649 => x"0266d47d",
   650 => x"66d487c7",
   651 => x"c505bf97",
   652 => x"c148c087",
   653 => x"66d487cf",
   654 => x"87f1fd49",
   655 => x"029c4c70",
   656 => x"dc87c0c1",
   657 => x"7d6949a4",
   658 => x"c449a4da",
   659 => x"699f4aa3",
   660 => x"d2c2c47a",
   661 => x"87d202bf",
   662 => x"9f49a4d4",
   663 => x"ffc04969",
   664 => x"487199ff",
   665 => x"7e7030d0",
   666 => x"7ec087c2",
   667 => x"6a48496e",
   668 => x"c07a7080",
   669 => x"49a3cc7b",
   670 => x"a3d0796a",
   671 => x"7479c049",
   672 => x"c087c248",
   673 => x"eafa2648",
   674 => x"5b5e0e87",
   675 => x"710e5d5c",
   676 => x"f1fec04c",
   677 => x"7478ff48",
   678 => x"cac1029c",
   679 => x"49a4c887",
   680 => x"c2c10269",
   681 => x"4a66d087",
   682 => x"d482496c",
   683 => x"66d05aa6",
   684 => x"c2c4b94d",
   685 => x"ff4abfce",
   686 => x"719972ba",
   687 => x"e4c00299",
   688 => x"4ba4c487",
   689 => x"f2f9496b",
   690 => x"c47b7087",
   691 => x"49bfcac2",
   692 => x"7c71816c",
   693 => x"c2c4b975",
   694 => x"ff4abfce",
   695 => x"719972ba",
   696 => x"dcff0599",
   697 => x"f97c7587",
   698 => x"731e87c9",
   699 => x"9b4b711e",
   700 => x"c887c702",
   701 => x"056949a3",
   702 => x"48c087c5",
   703 => x"c487ebc0",
   704 => x"4abfe3c6",
   705 => x"6949a3c4",
   706 => x"c489c249",
   707 => x"91bfcac2",
   708 => x"c44aa271",
   709 => x"49bfcec2",
   710 => x"a271996b",
   711 => x"1e66c84a",
   712 => x"d0ea4972",
   713 => x"7086c487",
   714 => x"caf84849",
   715 => x"1e731e87",
   716 => x"029b4b71",
   717 => x"a3c887c7",
   718 => x"c5056949",
   719 => x"c048c087",
   720 => x"c6c487eb",
   721 => x"c44abfe3",
   722 => x"496949a3",
   723 => x"c2c489c2",
   724 => x"7191bfca",
   725 => x"c2c44aa2",
   726 => x"6b49bfce",
   727 => x"4aa27199",
   728 => x"721e66c8",
   729 => x"87c3e649",
   730 => x"497086c4",
   731 => x"87c7f748",
   732 => x"5c5b5e0e",
   733 => x"711e0e5d",
   734 => x"4c66d44b",
   735 => x"9b732cc9",
   736 => x"87cfc102",
   737 => x"6949a3c8",
   738 => x"87c7c102",
   739 => x"d44da3d0",
   740 => x"c2c47d66",
   741 => x"ff49bfce",
   742 => x"994a6bb9",
   743 => x"03ac717e",
   744 => x"7bc087cd",
   745 => x"4aa3cc7d",
   746 => x"6a49a3c4",
   747 => x"7287c279",
   748 => x"029c748c",
   749 => x"1e4987dd",
   750 => x"ccfb4973",
   751 => x"d486c487",
   752 => x"ffc74966",
   753 => x"87cb0299",
   754 => x"1ecafac3",
   755 => x"d9fc4973",
   756 => x"2686c487",
   757 => x"0e87dcf5",
   758 => x"5d5c5b5e",
   759 => x"d086f00e",
   760 => x"e4c059a6",
   761 => x"66cc4b66",
   762 => x"4887ca02",
   763 => x"7e7080c8",
   764 => x"c505bf6e",
   765 => x"c348c087",
   766 => x"66cc87ec",
   767 => x"7384d04c",
   768 => x"48a6c449",
   769 => x"66c4786c",
   770 => x"6e80c481",
   771 => x"66c878bf",
   772 => x"87c606a9",
   773 => x"8966c449",
   774 => x"b7c04b71",
   775 => x"87c401ab",
   776 => x"87c2c348",
   777 => x"c74866c4",
   778 => x"7e7098ff",
   779 => x"c9c1026e",
   780 => x"49c0c887",
   781 => x"4a71896e",
   782 => x"4dcafac3",
   783 => x"b773856e",
   784 => x"87c106aa",
   785 => x"4849724a",
   786 => x"708066c4",
   787 => x"498b727c",
   788 => x"99718ac1",
   789 => x"c087d902",
   790 => x"154866e0",
   791 => x"66e0c050",
   792 => x"c080c148",
   793 => x"7258a6e4",
   794 => x"718ac149",
   795 => x"87e70599",
   796 => x"66d01ec1",
   797 => x"87d1f849",
   798 => x"b7c086c4",
   799 => x"e3c106ab",
   800 => x"66e0c087",
   801 => x"b7ffc74d",
   802 => x"e2c006ab",
   803 => x"d01e7587",
   804 => x"d5f94966",
   805 => x"85c0c887",
   806 => x"c0c8486c",
   807 => x"c87c7080",
   808 => x"1ec18bc0",
   809 => x"f74966d4",
   810 => x"86c887df",
   811 => x"c387eec0",
   812 => x"d01ecafa",
   813 => x"f1f84966",
   814 => x"c386c487",
   815 => x"734acafa",
   816 => x"806c4849",
   817 => x"49737c70",
   818 => x"99718bc1",
   819 => x"1287ce02",
   820 => x"85c17d97",
   821 => x"8bc14973",
   822 => x"f2059971",
   823 => x"abb7c087",
   824 => x"87e1fe01",
   825 => x"8ef048c1",
   826 => x"0e87c8f1",
   827 => x"5d5c5b5e",
   828 => x"9b4b710e",
   829 => x"c887c702",
   830 => x"056d4da3",
   831 => x"48ff87c5",
   832 => x"d087fdc0",
   833 => x"496c4ca3",
   834 => x"0599ffc7",
   835 => x"026c87d8",
   836 => x"1ec187c9",
   837 => x"f0f54973",
   838 => x"c386c487",
   839 => x"731ecafa",
   840 => x"87c6f749",
   841 => x"4a6c86c4",
   842 => x"c404aa6d",
   843 => x"cf48ff87",
   844 => x"7ca2c187",
   845 => x"ffc74972",
   846 => x"cafac399",
   847 => x"48699781",
   848 => x"1e87f0ef",
   849 => x"4b711e73",
   850 => x"e4c0029b",
   851 => x"f7c6c487",
   852 => x"c24a735b",
   853 => x"cac2c48a",
   854 => x"c49249bf",
   855 => x"48bfe3c6",
   856 => x"c6c48072",
   857 => x"487158fb",
   858 => x"c2c430c4",
   859 => x"edc058da",
   860 => x"f3c6c487",
   861 => x"e7c6c448",
   862 => x"c6c478bf",
   863 => x"c6c448f7",
   864 => x"c478bfeb",
   865 => x"02bfd2c2",
   866 => x"c2c487c9",
   867 => x"c449bfca",
   868 => x"c487c731",
   869 => x"49bfefc6",
   870 => x"c2c431c4",
   871 => x"d6ee59da",
   872 => x"5b5e0e87",
   873 => x"4a710e5c",
   874 => x"9a724bc0",
   875 => x"87e1c002",
   876 => x"9f49a2da",
   877 => x"c2c44b69",
   878 => x"cf02bfd2",
   879 => x"49a2d487",
   880 => x"4c49699f",
   881 => x"9cffffc0",
   882 => x"87c234d0",
   883 => x"49744cc0",
   884 => x"fd4973b3",
   885 => x"dced87ed",
   886 => x"5b5e0e87",
   887 => x"f40e5d5c",
   888 => x"c04a7186",
   889 => x"029a727e",
   890 => x"fac387d8",
   891 => x"78c048c6",
   892 => x"48fef9c3",
   893 => x"bff7c6c4",
   894 => x"c2fac378",
   895 => x"f3c6c448",
   896 => x"c2c478bf",
   897 => x"50c048e7",
   898 => x"bfd6c2c4",
   899 => x"c6fac349",
   900 => x"aa714abf",
   901 => x"87c0c403",
   902 => x"99cf4972",
   903 => x"87e1c005",
   904 => x"1ecafac3",
   905 => x"bffef9c3",
   906 => x"fef9c349",
   907 => x"78a1c148",
   908 => x"c0deff71",
   909 => x"c086c487",
   910 => x"c348edfe",
   911 => x"cc78cafa",
   912 => x"edfec087",
   913 => x"e0c048bf",
   914 => x"f1fec080",
   915 => x"c6fac358",
   916 => x"80c148bf",
   917 => x"58cafac3",
   918 => x"000fad27",
   919 => x"bf97bf00",
   920 => x"c2029d4d",
   921 => x"e5c387e2",
   922 => x"dbc202ad",
   923 => x"edfec087",
   924 => x"a3cb4bbf",
   925 => x"cf4c1149",
   926 => x"d2c105ac",
   927 => x"df497587",
   928 => x"cd89c199",
   929 => x"dac2c491",
   930 => x"4aa3c181",
   931 => x"a3c35112",
   932 => x"c551124a",
   933 => x"51124aa3",
   934 => x"124aa3c7",
   935 => x"4aa3c951",
   936 => x"a3ce5112",
   937 => x"d051124a",
   938 => x"51124aa3",
   939 => x"124aa3d2",
   940 => x"4aa3d451",
   941 => x"a3d65112",
   942 => x"d851124a",
   943 => x"51124aa3",
   944 => x"124aa3dc",
   945 => x"4aa3de51",
   946 => x"7ec15112",
   947 => x"7487f9c0",
   948 => x"0599c849",
   949 => x"7487eac0",
   950 => x"0599d049",
   951 => x"66dc87d0",
   952 => x"87cac002",
   953 => x"66dc4973",
   954 => x"0298700f",
   955 => x"056e87d3",
   956 => x"c487c6c0",
   957 => x"c048dac2",
   958 => x"edfec050",
   959 => x"e7c248bf",
   960 => x"e7c2c487",
   961 => x"7e50c048",
   962 => x"bfd6c2c4",
   963 => x"c6fac349",
   964 => x"aa714abf",
   965 => x"87c0fc04",
   966 => x"bff7c6c4",
   967 => x"87c8c005",
   968 => x"bfd2c2c4",
   969 => x"87fec102",
   970 => x"48f1fec0",
   971 => x"fac378ff",
   972 => x"e849bfc2",
   973 => x"497087c5",
   974 => x"59c6fac3",
   975 => x"c348a6c4",
   976 => x"78bfc2fa",
   977 => x"bfd2c2c4",
   978 => x"87d8c002",
   979 => x"cf4966c4",
   980 => x"f8ffffff",
   981 => x"c002a999",
   982 => x"4dc087c5",
   983 => x"c187e1c0",
   984 => x"87dcc04d",
   985 => x"cf4966c4",
   986 => x"a999f8ff",
   987 => x"87c8c002",
   988 => x"c048a6c8",
   989 => x"87c5c078",
   990 => x"c148a6c8",
   991 => x"4d66c878",
   992 => x"c0059d75",
   993 => x"66c487e0",
   994 => x"c489c249",
   995 => x"4abfcac2",
   996 => x"e3c6c491",
   997 => x"f9c34abf",
   998 => x"a17248fe",
   999 => x"c6fac378",
  1000 => x"f978c048",
  1001 => x"48c087e2",
  1002 => x"c6e68ef4",
  1003 => x"00000087",
  1004 => x"ffffff00",
  1005 => x"000fbdff",
  1006 => x"000fc600",
  1007 => x"54414600",
  1008 => x"20203233",
  1009 => x"41460020",
  1010 => x"20363154",
  1011 => x"1e002020",
  1012 => x"c348d4ff",
  1013 => x"486878ff",
  1014 => x"ff1e4f26",
  1015 => x"ffc348d4",
  1016 => x"48d0ff78",
  1017 => x"ff78e1c8",
  1018 => x"78d448d4",
  1019 => x"48fbc6c4",
  1020 => x"50bfd4ff",
  1021 => x"ff1e4f26",
  1022 => x"e0c048d0",
  1023 => x"1e4f2678",
  1024 => x"7087ccff",
  1025 => x"c6029949",
  1026 => x"a9fbc087",
  1027 => x"7187f105",
  1028 => x"0e4f2648",
  1029 => x"0e5c5b5e",
  1030 => x"4cc04b71",
  1031 => x"7087f0fe",
  1032 => x"c0029949",
  1033 => x"ecc087f9",
  1034 => x"f2c002a9",
  1035 => x"a9fbc087",
  1036 => x"87ebc002",
  1037 => x"acb766cc",
  1038 => x"d087c703",
  1039 => x"87c20266",
  1040 => x"99715371",
  1041 => x"c187c202",
  1042 => x"87c3fe84",
  1043 => x"02994970",
  1044 => x"ecc087cd",
  1045 => x"87c702a9",
  1046 => x"05a9fbc0",
  1047 => x"d087d5ff",
  1048 => x"87c30266",
  1049 => x"c07b97c0",
  1050 => x"c405a9ec",
  1051 => x"c54a7487",
  1052 => x"c04a7487",
  1053 => x"48728a0a",
  1054 => x"4d2687c2",
  1055 => x"4b264c26",
  1056 => x"fd1e4f26",
  1057 => x"497087c9",
  1058 => x"a9b7f0c0",
  1059 => x"c087ca04",
  1060 => x"01a9b7f9",
  1061 => x"f0c087c3",
  1062 => x"b7c1c189",
  1063 => x"87ca04a9",
  1064 => x"a9b7dac1",
  1065 => x"c087c301",
  1066 => x"487189f7",
  1067 => x"5e0e4f26",
  1068 => x"710e5c5b",
  1069 => x"4cd4ff4a",
  1070 => x"eac04972",
  1071 => x"9b4b7087",
  1072 => x"c187c202",
  1073 => x"48d0ff8b",
  1074 => x"c178c5c8",
  1075 => x"49737cd5",
  1076 => x"f7c331c6",
  1077 => x"4abf97fc",
  1078 => x"70b07148",
  1079 => x"48d0ff7c",
  1080 => x"487378c4",
  1081 => x"0e87d5fe",
  1082 => x"5d5c5b5e",
  1083 => x"7186f80e",
  1084 => x"fb7ec04c",
  1085 => x"4bc087e4",
  1086 => x"97d4c6c1",
  1087 => x"a9c049bf",
  1088 => x"fb87cf04",
  1089 => x"83c187f9",
  1090 => x"97d4c6c1",
  1091 => x"06ab49bf",
  1092 => x"c6c187f1",
  1093 => x"02bf97d4",
  1094 => x"f2fa87cf",
  1095 => x"99497087",
  1096 => x"c087c602",
  1097 => x"f105a9ec",
  1098 => x"fa4bc087",
  1099 => x"4d7087e1",
  1100 => x"c887dcfa",
  1101 => x"d6fa58a6",
  1102 => x"c14a7087",
  1103 => x"49a4c883",
  1104 => x"ad496997",
  1105 => x"c087c702",
  1106 => x"c005adff",
  1107 => x"a4c987e7",
  1108 => x"49699749",
  1109 => x"02a966c4",
  1110 => x"c04887c7",
  1111 => x"d405a8ff",
  1112 => x"49a4ca87",
  1113 => x"aa496997",
  1114 => x"c087c602",
  1115 => x"c405aaff",
  1116 => x"d07ec187",
  1117 => x"adecc087",
  1118 => x"c087c602",
  1119 => x"c405adfb",
  1120 => x"c14bc087",
  1121 => x"fe026e7e",
  1122 => x"e9f987e1",
  1123 => x"f8487387",
  1124 => x"87e6fb8e",
  1125 => x"5b5e0e00",
  1126 => x"1e0e5d5c",
  1127 => x"4cc04b71",
  1128 => x"c004ab4d",
  1129 => x"c3c187e8",
  1130 => x"9d751ee7",
  1131 => x"c087c402",
  1132 => x"c187c24a",
  1133 => x"f049724a",
  1134 => x"86c487df",
  1135 => x"84c17e70",
  1136 => x"87c2056e",
  1137 => x"85c14c73",
  1138 => x"ff06ac73",
  1139 => x"486e87d8",
  1140 => x"264d2626",
  1141 => x"264b264c",
  1142 => x"4a711e4f",
  1143 => x"99ffc349",
  1144 => x"7148d4ff",
  1145 => x"c8497278",
  1146 => x"ffc329b7",
  1147 => x"72787199",
  1148 => x"29b7d049",
  1149 => x"7199ffc3",
  1150 => x"d8497278",
  1151 => x"ffc329b7",
  1152 => x"26787199",
  1153 => x"5b5e0e4f",
  1154 => x"1e0e5d5c",
  1155 => x"4bc04a71",
  1156 => x"e3c14972",
  1157 => x"987087d6",
  1158 => x"c187da05",
  1159 => x"c149744c",
  1160 => x"7087e3e4",
  1161 => x"87c20598",
  1162 => x"84c14bc1",
  1163 => x"bfdecbc4",
  1164 => x"e806acb7",
  1165 => x"48d0ff87",
  1166 => x"ff78e1c8",
  1167 => x"78dd48d4",
  1168 => x"c7029b73",
  1169 => x"c6ccc487",
  1170 => x"87c24dbf",
  1171 => x"49754dc0",
  1172 => x"7387c6fe",
  1173 => x"87c7029b",
  1174 => x"bfc6ccc4",
  1175 => x"c087c27e",
  1176 => x"fd496e7e",
  1177 => x"49c087f3",
  1178 => x"c087eefd",
  1179 => x"87e9fd49",
  1180 => x"c048d0ff",
  1181 => x"1ec178e0",
  1182 => x"f2c049dc",
  1183 => x"487387db",
  1184 => x"ccfd8ef8",
  1185 => x"5b5e0e87",
  1186 => x"1e0e5d5c",
  1187 => x"de494c71",
  1188 => x"d5c7c491",
  1189 => x"9785714d",
  1190 => x"ddc1026d",
  1191 => x"c0c7c487",
  1192 => x"82744abf",
  1193 => x"ecfb4972",
  1194 => x"6e7e7087",
  1195 => x"87f3c002",
  1196 => x"4bc8c7c4",
  1197 => x"49cb4a6e",
  1198 => x"87fdf7fe",
  1199 => x"93cb4b74",
  1200 => x"83e4edc1",
  1201 => x"cbc183c4",
  1202 => x"49747bfe",
  1203 => x"87ffc4c1",
  1204 => x"c7c47b75",
  1205 => x"49bf97d4",
  1206 => x"c8c7c41e",
  1207 => x"d0ebc249",
  1208 => x"7486c487",
  1209 => x"e6c4c149",
  1210 => x"c149c087",
  1211 => x"c487c5c6",
  1212 => x"c048fcc6",
  1213 => x"dd49c178",
  1214 => x"fb2687d2",
  1215 => x"6f4c87d3",
  1216 => x"6e696461",
  1217 => x"2e2e2e67",
  1218 => x"5b5e0e00",
  1219 => x"4b710e5c",
  1220 => x"c0c7c44a",
  1221 => x"497282bf",
  1222 => x"7087faf9",
  1223 => x"c4029c4c",
  1224 => x"fce94987",
  1225 => x"c0c7c487",
  1226 => x"c178c048",
  1227 => x"87dcdc49",
  1228 => x"0e87e0fa",
  1229 => x"5d5c5b5e",
  1230 => x"c386f40e",
  1231 => x"c04dcafa",
  1232 => x"48a6c44c",
  1233 => x"c7c478c0",
  1234 => x"c049bfc0",
  1235 => x"c1c106a9",
  1236 => x"cafac387",
  1237 => x"c0029848",
  1238 => x"c3c187f8",
  1239 => x"66c81ee7",
  1240 => x"c487c702",
  1241 => x"78c048a6",
  1242 => x"a6c487c5",
  1243 => x"c478c148",
  1244 => x"e4e94966",
  1245 => x"7086c487",
  1246 => x"c484c14d",
  1247 => x"80c14866",
  1248 => x"c458a6c8",
  1249 => x"49bfc0c7",
  1250 => x"87c603ac",
  1251 => x"ff059d75",
  1252 => x"4cc087c8",
  1253 => x"c3029d75",
  1254 => x"c3c187e0",
  1255 => x"66c81ee7",
  1256 => x"cc87c702",
  1257 => x"78c048a6",
  1258 => x"a6cc87c5",
  1259 => x"cc78c148",
  1260 => x"e4e84966",
  1261 => x"7086c487",
  1262 => x"c2026e7e",
  1263 => x"496e87e9",
  1264 => x"699781cb",
  1265 => x"0299d049",
  1266 => x"c187d6c1",
  1267 => x"744ac9cc",
  1268 => x"c191cb49",
  1269 => x"7281e4ed",
  1270 => x"c381c879",
  1271 => x"497451ff",
  1272 => x"c7c491de",
  1273 => x"85714dd5",
  1274 => x"7d97c1c2",
  1275 => x"c049a5c1",
  1276 => x"c2c451e0",
  1277 => x"02bf97da",
  1278 => x"84c187d2",
  1279 => x"c44ba5c2",
  1280 => x"db4adac2",
  1281 => x"f0f2fe49",
  1282 => x"87dbc187",
  1283 => x"c049a5cd",
  1284 => x"c284c151",
  1285 => x"4a6e4ba5",
  1286 => x"f2fe49cb",
  1287 => x"c6c187db",
  1288 => x"c5cac187",
  1289 => x"cb49744a",
  1290 => x"e4edc191",
  1291 => x"c4797281",
  1292 => x"bf97dac2",
  1293 => x"7487d802",
  1294 => x"c191de49",
  1295 => x"d5c7c484",
  1296 => x"c483714b",
  1297 => x"dd4adac2",
  1298 => x"ecf1fe49",
  1299 => x"7487d887",
  1300 => x"c493de4b",
  1301 => x"cb83d5c7",
  1302 => x"51c049a3",
  1303 => x"6e7384c1",
  1304 => x"fe49cb4a",
  1305 => x"c487d2f1",
  1306 => x"80c14866",
  1307 => x"c758a6c8",
  1308 => x"c5c003ac",
  1309 => x"fc056e87",
  1310 => x"487487e0",
  1311 => x"d0f58ef4",
  1312 => x"1e731e87",
  1313 => x"cb494b71",
  1314 => x"e4edc191",
  1315 => x"4aa1c881",
  1316 => x"48fcf7c3",
  1317 => x"a1c95012",
  1318 => x"d4c6c14a",
  1319 => x"ca501248",
  1320 => x"d4c7c481",
  1321 => x"c4501148",
  1322 => x"bf97d4c7",
  1323 => x"49c01e49",
  1324 => x"87fde3c2",
  1325 => x"48fcc6c4",
  1326 => x"49c178de",
  1327 => x"2687cdd6",
  1328 => x"1e87d2f4",
  1329 => x"cb494a71",
  1330 => x"e4edc191",
  1331 => x"1181c881",
  1332 => x"c0c7c448",
  1333 => x"c0c7c458",
  1334 => x"c178c048",
  1335 => x"87ecd549",
  1336 => x"c01e4f26",
  1337 => x"cbfec049",
  1338 => x"1e4f2687",
  1339 => x"d2029971",
  1340 => x"f9eec187",
  1341 => x"f750c048",
  1342 => x"c3d3c180",
  1343 => x"ddedc140",
  1344 => x"c187ce78",
  1345 => x"c148f5ee",
  1346 => x"fc78d6ed",
  1347 => x"e2d3c180",
  1348 => x"0e4f2678",
  1349 => x"0e5c5b5e",
  1350 => x"cb4a4c71",
  1351 => x"e4edc192",
  1352 => x"49a2c882",
  1353 => x"974ba2c9",
  1354 => x"971e4b6b",
  1355 => x"ca1e4969",
  1356 => x"c0491282",
  1357 => x"c087c6e9",
  1358 => x"87d0d449",
  1359 => x"fbc04974",
  1360 => x"8ef887cd",
  1361 => x"1e87ccf2",
  1362 => x"4b711e73",
  1363 => x"87c3ff49",
  1364 => x"fefe4973",
  1365 => x"87fdf187",
  1366 => x"711e731e",
  1367 => x"4aa3c64b",
  1368 => x"c187db02",
  1369 => x"87d6028a",
  1370 => x"dac1028a",
  1371 => x"c0028a87",
  1372 => x"028a87fc",
  1373 => x"8a87e1c0",
  1374 => x"c187cb02",
  1375 => x"49c787db",
  1376 => x"c187c0fd",
  1377 => x"c7c487de",
  1378 => x"c102bfc0",
  1379 => x"c14887cb",
  1380 => x"c4c7c488",
  1381 => x"87c1c158",
  1382 => x"bfc4c7c4",
  1383 => x"87f9c002",
  1384 => x"bfc0c7c4",
  1385 => x"c480c148",
  1386 => x"c058c4c7",
  1387 => x"c7c487eb",
  1388 => x"c649bfc0",
  1389 => x"c4c7c489",
  1390 => x"a9b7c059",
  1391 => x"c487da03",
  1392 => x"c048c0c7",
  1393 => x"c487d278",
  1394 => x"02bfc4c7",
  1395 => x"c7c487cb",
  1396 => x"c648bfc0",
  1397 => x"c4c7c480",
  1398 => x"d149c058",
  1399 => x"497387ee",
  1400 => x"87ebf8c0",
  1401 => x"0e87eeef",
  1402 => x"0e5c5b5e",
  1403 => x"66cc4c71",
  1404 => x"cb4b741e",
  1405 => x"e4edc193",
  1406 => x"4aa3c483",
  1407 => x"ebfe496a",
  1408 => x"d2c187c7",
  1409 => x"a3c87bc1",
  1410 => x"5166d449",
  1411 => x"d849a3c9",
  1412 => x"a3ca5166",
  1413 => x"5166dc49",
  1414 => x"87f7ee26",
  1415 => x"5c5b5e0e",
  1416 => x"d0ff0e5d",
  1417 => x"59a6d886",
  1418 => x"c048a6c4",
  1419 => x"c180c478",
  1420 => x"c47866c4",
  1421 => x"c478c180",
  1422 => x"c478c180",
  1423 => x"c148c4c7",
  1424 => x"fcc6c478",
  1425 => x"a8de48bf",
  1426 => x"f387cb05",
  1427 => x"497087e5",
  1428 => x"ce59a6c8",
  1429 => x"c1e687fe",
  1430 => x"87e3e687",
  1431 => x"7087f0e5",
  1432 => x"acfbc04c",
  1433 => x"87d0c102",
  1434 => x"c10566d4",
  1435 => x"1ec087c2",
  1436 => x"c11ec11e",
  1437 => x"c01ed7ef",
  1438 => x"87ebfd49",
  1439 => x"4a66d0c1",
  1440 => x"496a82c4",
  1441 => x"517481c7",
  1442 => x"1ed81ec1",
  1443 => x"81c8496a",
  1444 => x"d887c0e6",
  1445 => x"66c4c186",
  1446 => x"01a8c048",
  1447 => x"a6c487c7",
  1448 => x"ce78c148",
  1449 => x"66c4c187",
  1450 => x"cc88c148",
  1451 => x"87c358a6",
  1452 => x"cc87cce5",
  1453 => x"78c248a6",
  1454 => x"cd029c74",
  1455 => x"66c487d2",
  1456 => x"66c8c148",
  1457 => x"c7cd03a8",
  1458 => x"48a6d887",
  1459 => x"fee378c0",
  1460 => x"c14c7087",
  1461 => x"c205acd0",
  1462 => x"66d887d6",
  1463 => x"87e2e67e",
  1464 => x"a6dc4970",
  1465 => x"87e7e359",
  1466 => x"ecc04c70",
  1467 => x"eac105ac",
  1468 => x"4966c487",
  1469 => x"c0c191cb",
  1470 => x"a1c48166",
  1471 => x"c84d6a4a",
  1472 => x"66d84aa1",
  1473 => x"c3d3c152",
  1474 => x"87c3e379",
  1475 => x"029c4c70",
  1476 => x"fbc087d8",
  1477 => x"87d202ac",
  1478 => x"f2e25574",
  1479 => x"9c4c7087",
  1480 => x"c087c702",
  1481 => x"ff05acfb",
  1482 => x"e0c087ee",
  1483 => x"55c1c255",
  1484 => x"d47d97c0",
  1485 => x"a96e4966",
  1486 => x"c487db05",
  1487 => x"66c84866",
  1488 => x"87ca04a8",
  1489 => x"c14866c4",
  1490 => x"58a6c880",
  1491 => x"66c887c8",
  1492 => x"cc88c148",
  1493 => x"f6e158a6",
  1494 => x"c14c7087",
  1495 => x"c805acd0",
  1496 => x"4866d087",
  1497 => x"a6d480c1",
  1498 => x"acd0c158",
  1499 => x"87eafd02",
  1500 => x"d448a6dc",
  1501 => x"66d87866",
  1502 => x"a866dc48",
  1503 => x"87e2c905",
  1504 => x"48a6e0c0",
  1505 => x"c478f0c0",
  1506 => x"7866cc80",
  1507 => x"78c080c4",
  1508 => x"c048747e",
  1509 => x"f0c088fb",
  1510 => x"987058a6",
  1511 => x"87ddc802",
  1512 => x"c088cb48",
  1513 => x"7058a6f0",
  1514 => x"e9c00298",
  1515 => x"88c94887",
  1516 => x"58a6f0c0",
  1517 => x"c3029870",
  1518 => x"c44887e5",
  1519 => x"a6f0c088",
  1520 => x"02987058",
  1521 => x"c14887de",
  1522 => x"a6f0c088",
  1523 => x"02987058",
  1524 => x"c787ccc3",
  1525 => x"e0c087e1",
  1526 => x"78c048a6",
  1527 => x"c14866cc",
  1528 => x"58a6d080",
  1529 => x"87e7dfff",
  1530 => x"ecc04c70",
  1531 => x"87d502ac",
  1532 => x"0266e0c0",
  1533 => x"e4c087c6",
  1534 => x"87c95ca6",
  1535 => x"f0c04874",
  1536 => x"a6e8c088",
  1537 => x"acecc058",
  1538 => x"ff87cd02",
  1539 => x"7087c0df",
  1540 => x"acecc04c",
  1541 => x"87f3ff05",
  1542 => x"1e66e0c0",
  1543 => x"1e4966d4",
  1544 => x"1e66ecc0",
  1545 => x"1ed7efc1",
  1546 => x"f64966d4",
  1547 => x"1ec087f9",
  1548 => x"66dc1eca",
  1549 => x"c191cb49",
  1550 => x"d88166d8",
  1551 => x"a1c448a6",
  1552 => x"bf66d878",
  1553 => x"cadfff49",
  1554 => x"c086d887",
  1555 => x"c106a8b7",
  1556 => x"1ec187c8",
  1557 => x"66c81ede",
  1558 => x"deff49bf",
  1559 => x"86c887f5",
  1560 => x"c0484970",
  1561 => x"e4c08808",
  1562 => x"b7c058a6",
  1563 => x"e9c006a8",
  1564 => x"66e0c087",
  1565 => x"a8b7dd48",
  1566 => x"6e87df03",
  1567 => x"e0c049bf",
  1568 => x"e0c08166",
  1569 => x"c1496651",
  1570 => x"81bf6e81",
  1571 => x"c051c1c2",
  1572 => x"c24966e0",
  1573 => x"81bf6e81",
  1574 => x"7ec151c0",
  1575 => x"ff87dec4",
  1576 => x"c087dfdf",
  1577 => x"ff58a6e4",
  1578 => x"c087d7df",
  1579 => x"c058a6e8",
  1580 => x"c005a8ec",
  1581 => x"e4c087cb",
  1582 => x"e0c048a6",
  1583 => x"c4c07866",
  1584 => x"cadcff87",
  1585 => x"4966c487",
  1586 => x"c0c191cb",
  1587 => x"80714866",
  1588 => x"4a6e7e70",
  1589 => x"496e82c8",
  1590 => x"e0c081ca",
  1591 => x"e4c05166",
  1592 => x"81c14966",
  1593 => x"8966e0c0",
  1594 => x"307148c1",
  1595 => x"89c14970",
  1596 => x"c47a9771",
  1597 => x"49bff1ca",
  1598 => x"2966e0c0",
  1599 => x"484a6a97",
  1600 => x"f0c09871",
  1601 => x"496e58a6",
  1602 => x"4d6981c4",
  1603 => x"d84866dc",
  1604 => x"c002a866",
  1605 => x"a6d887c8",
  1606 => x"c078c048",
  1607 => x"a6d887c5",
  1608 => x"d878c148",
  1609 => x"e0c01e66",
  1610 => x"ff49751e",
  1611 => x"c887e4db",
  1612 => x"c04c7086",
  1613 => x"c106acb7",
  1614 => x"857487d4",
  1615 => x"7449e0c0",
  1616 => x"c14b7589",
  1617 => x"714ac9e9",
  1618 => x"87edddfe",
  1619 => x"e8c085c2",
  1620 => x"80c14866",
  1621 => x"58a6ecc0",
  1622 => x"4966ecc0",
  1623 => x"a97081c1",
  1624 => x"87c8c002",
  1625 => x"c048a6d8",
  1626 => x"87c5c078",
  1627 => x"c148a6d8",
  1628 => x"1e66d878",
  1629 => x"c049a4c2",
  1630 => x"887148e0",
  1631 => x"751e4970",
  1632 => x"cedaff49",
  1633 => x"c086c887",
  1634 => x"ff01a8b7",
  1635 => x"e8c087c0",
  1636 => x"d1c00266",
  1637 => x"c9496e87",
  1638 => x"66e8c081",
  1639 => x"c1486e51",
  1640 => x"c078d3d4",
  1641 => x"496e87cc",
  1642 => x"51c281c9",
  1643 => x"d5c1486e",
  1644 => x"7ec178c7",
  1645 => x"ff87c6c0",
  1646 => x"7087c4d9",
  1647 => x"c0026e4c",
  1648 => x"66c487f5",
  1649 => x"a866c848",
  1650 => x"87cbc004",
  1651 => x"c14866c4",
  1652 => x"58a6c880",
  1653 => x"c887e0c0",
  1654 => x"88c14866",
  1655 => x"c058a6cc",
  1656 => x"c6c187d5",
  1657 => x"c8c005ac",
  1658 => x"4866cc87",
  1659 => x"a6d080c1",
  1660 => x"cad8ff58",
  1661 => x"d04c7087",
  1662 => x"80c14866",
  1663 => x"7458a6d4",
  1664 => x"cbc0029c",
  1665 => x"4866c487",
  1666 => x"a866c8c1",
  1667 => x"87f9f204",
  1668 => x"87e2d7ff",
  1669 => x"c74866c4",
  1670 => x"e5c003a8",
  1671 => x"c4c7c487",
  1672 => x"c478c048",
  1673 => x"91cb4966",
  1674 => x"8166c0c1",
  1675 => x"6a4aa1c4",
  1676 => x"7952c04a",
  1677 => x"c14866c4",
  1678 => x"58a6c880",
  1679 => x"ff04a8c7",
  1680 => x"d0ff87db",
  1681 => x"c8deff8e",
  1682 => x"00203a87",
  1683 => x"711e731e",
  1684 => x"c6029b4b",
  1685 => x"c0c7c487",
  1686 => x"c778c048",
  1687 => x"c0c7c41e",
  1688 => x"c11e49bf",
  1689 => x"c41ee4ed",
  1690 => x"49bffcc6",
  1691 => x"cc87edee",
  1692 => x"fcc6c486",
  1693 => x"f2e949bf",
  1694 => x"029b7387",
  1695 => x"edc187c8",
  1696 => x"e7c049e4",
  1697 => x"ddff87db",
  1698 => x"731e87cb",
  1699 => x"c34bc01e",
  1700 => x"c048fcf7",
  1701 => x"c7efc150",
  1702 => x"c8c249bf",
  1703 => x"987087e6",
  1704 => x"c187c405",
  1705 => x"734bedea",
  1706 => x"e8dcff48",
  1707 => x"4d4f5287",
  1708 => x"616f6c20",
  1709 => x"676e6964",
  1710 => x"69616620",
  1711 => x"0064656c",
  1712 => x"87f2c71e",
  1713 => x"c3fe49c1",
  1714 => x"ede6fe87",
  1715 => x"02987087",
  1716 => x"effe87cd",
  1717 => x"987087ea",
  1718 => x"c187c402",
  1719 => x"c087c24a",
  1720 => x"059a724a",
  1721 => x"1ec087ce",
  1722 => x"49d4ecc1",
  1723 => x"87c1f3c0",
  1724 => x"87fe86c4",
  1725 => x"87eeccc2",
  1726 => x"ecc11ec0",
  1727 => x"f2c049df",
  1728 => x"1ec087ef",
  1729 => x"7087c3fe",
  1730 => x"e4f2c049",
  1731 => x"87e5c387",
  1732 => x"4f268ef8",
  1733 => x"66204453",
  1734 => x"656c6961",
  1735 => x"42002e64",
  1736 => x"69746f6f",
  1737 => x"2e2e676e",
  1738 => x"c11e002e",
  1739 => x"c087c2fc",
  1740 => x"c187cce9",
  1741 => x"c287fafb",
  1742 => x"ee87f8c0",
  1743 => x"1e4f2687",
  1744 => x"48c0c7c4",
  1745 => x"c6c478c0",
  1746 => x"78c048fc",
  1747 => x"ff87f1fd",
  1748 => x"48c087d8",
  1749 => x"20804f26",
  1750 => x"74697845",
  1751 => x"42208000",
  1752 => x"006b6361",
  1753 => x"000014c3",
  1754 => x"000041d5",
  1755 => x"c3000000",
  1756 => x"f3000014",
  1757 => x"00000041",
  1758 => x"14c30000",
  1759 => x"42110000",
  1760 => x"00000000",
  1761 => x"0014c300",
  1762 => x"00422f00",
  1763 => x"00000000",
  1764 => x"000014c3",
  1765 => x"0000424d",
  1766 => x"c3000000",
  1767 => x"6b000014",
  1768 => x"00000042",
  1769 => x"14c30000",
  1770 => x"42890000",
  1771 => x"00000000",
  1772 => x"0014c300",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00001558",
  1776 => x"00000000",
  1777 => x"cb000000",
  1778 => x"4e00001b",
  1779 => x"45474f45",
  1780 => x"5220204f",
  1781 => x"4c004d4f",
  1782 => x"2064616f",
  1783 => x"1e002e2a",
  1784 => x"c048f0fe",
  1785 => x"7909cd78",
  1786 => x"1e4f2609",
  1787 => x"bff0fe1e",
  1788 => x"2626487e",
  1789 => x"f0fe1e4f",
  1790 => x"2678c148",
  1791 => x"f0fe1e4f",
  1792 => x"2678c048",
  1793 => x"4a711e4f",
  1794 => x"265252c0",
  1795 => x"5b5e0e4f",
  1796 => x"f40e5d5c",
  1797 => x"974d7186",
  1798 => x"a5c17e6d",
  1799 => x"486c974c",
  1800 => x"6e58a6c8",
  1801 => x"a866c448",
  1802 => x"ff87c505",
  1803 => x"87e6c048",
  1804 => x"c287caff",
  1805 => x"6c9749a5",
  1806 => x"4ba3714b",
  1807 => x"974b6b97",
  1808 => x"486e7e6c",
  1809 => x"a6c880c1",
  1810 => x"cc98c758",
  1811 => x"977058a6",
  1812 => x"87e1fe7c",
  1813 => x"8ef44873",
  1814 => x"4c264d26",
  1815 => x"4f264b26",
  1816 => x"5c5b5e0e",
  1817 => x"7186f40e",
  1818 => x"4a66d84c",
  1819 => x"c29affc3",
  1820 => x"6c974ba4",
  1821 => x"49a17349",
  1822 => x"6c975172",
  1823 => x"c1486e7e",
  1824 => x"58a6c880",
  1825 => x"a6cc98c7",
  1826 => x"f4547058",
  1827 => x"87caff8e",
  1828 => x"e8fd1e1e",
  1829 => x"4abfe087",
  1830 => x"c0e0c049",
  1831 => x"87cb0299",
  1832 => x"cac41e72",
  1833 => x"f7fe49e7",
  1834 => x"fc86c487",
  1835 => x"7e7087fd",
  1836 => x"2687c2fd",
  1837 => x"c41e4f26",
  1838 => x"fd49e7ca",
  1839 => x"f2c187c7",
  1840 => x"dafc49d0",
  1841 => x"87d5c687",
  1842 => x"5e0e4f26",
  1843 => x"0e5d5c5b",
  1844 => x"bfc6cbc4",
  1845 => x"def4c14a",
  1846 => x"724c49bf",
  1847 => x"fc4d71bc",
  1848 => x"4bc087db",
  1849 => x"99d04974",
  1850 => x"7587d502",
  1851 => x"7199d049",
  1852 => x"c11ec01e",
  1853 => x"734aecfb",
  1854 => x"c1491282",
  1855 => x"86c887ca",
  1856 => x"832d2cc1",
  1857 => x"ff04abc8",
  1858 => x"e8fb87da",
  1859 => x"def4c187",
  1860 => x"c6cbc448",
  1861 => x"4d2678bf",
  1862 => x"4b264c26",
  1863 => x"00004f26",
  1864 => x"731e0000",
  1865 => x"c04b711e",
  1866 => x"ecfbc14a",
  1867 => x"97817249",
  1868 => x"a9734969",
  1869 => x"c187c405",
  1870 => x"c187ca48",
  1871 => x"aab7c882",
  1872 => x"c087e604",
  1873 => x"87d2ff48",
  1874 => x"711e731e",
  1875 => x"d1ff494b",
  1876 => x"02987087",
  1877 => x"ff87ecc0",
  1878 => x"e1c848d0",
  1879 => x"48d4ff78",
  1880 => x"66c878c5",
  1881 => x"c387c302",
  1882 => x"66cc78e0",
  1883 => x"ff87c602",
  1884 => x"f0c348d4",
  1885 => x"48d4ff78",
  1886 => x"d0ff7873",
  1887 => x"78e1c848",
  1888 => x"fe78e0c0",
  1889 => x"5e0e87d4",
  1890 => x"710e5c5b",
  1891 => x"e7cac44c",
  1892 => x"87f9f949",
  1893 => x"b7c04a70",
  1894 => x"e3c204aa",
  1895 => x"aae0c387",
  1896 => x"c187c905",
  1897 => x"c148c9f9",
  1898 => x"87d4c278",
  1899 => x"05aaf0c3",
  1900 => x"f9c187c9",
  1901 => x"78c148c5",
  1902 => x"c187f5c1",
  1903 => x"02bfc9f9",
  1904 => x"4b7287c7",
  1905 => x"c2b3c0c2",
  1906 => x"744b7287",
  1907 => x"87d1059c",
  1908 => x"bfc5f9c1",
  1909 => x"c9f9c11e",
  1910 => x"49721ebf",
  1911 => x"c887e9fd",
  1912 => x"c5f9c186",
  1913 => x"e0c002bf",
  1914 => x"c4497387",
  1915 => x"c19129b7",
  1916 => x"7381ecfa",
  1917 => x"c29acf4a",
  1918 => x"7248c192",
  1919 => x"ff4a7030",
  1920 => x"694872ba",
  1921 => x"db797098",
  1922 => x"c4497387",
  1923 => x"c19129b7",
  1924 => x"7381ecfa",
  1925 => x"c29acf4a",
  1926 => x"7248c392",
  1927 => x"484a7030",
  1928 => x"7970b069",
  1929 => x"48c9f9c1",
  1930 => x"f9c178c0",
  1931 => x"78c048c5",
  1932 => x"49e7cac4",
  1933 => x"7087d6f7",
  1934 => x"aab7c04a",
  1935 => x"87ddfd03",
  1936 => x"d3fb48c0",
  1937 => x"00000087",
  1938 => x"00000000",
  1939 => x"1e731e00",
  1940 => x"f5f94b71",
  1941 => x"fc497387",
  1942 => x"fdfa87ec",
  1943 => x"4ac01e87",
  1944 => x"91c44972",
  1945 => x"81ecfac1",
  1946 => x"82c179c0",
  1947 => x"04aab7d0",
  1948 => x"4f2687ee",
  1949 => x"5c5b5e0e",
  1950 => x"4d710e5d",
  1951 => x"7587fef5",
  1952 => x"2ab7c44a",
  1953 => x"ecfac192",
  1954 => x"cf4c7582",
  1955 => x"6a94c29c",
  1956 => x"2b744b49",
  1957 => x"48c29bc3",
  1958 => x"4c703074",
  1959 => x"4874bcff",
  1960 => x"7a709871",
  1961 => x"7387cef5",
  1962 => x"87eaf948",
  1963 => x"00000000",
  1964 => x"00000000",
  1965 => x"00000000",
  1966 => x"00000000",
  1967 => x"00000000",
  1968 => x"00000000",
  1969 => x"00000000",
  1970 => x"00000000",
  1971 => x"00000000",
  1972 => x"00000000",
  1973 => x"00000000",
  1974 => x"00000000",
  1975 => x"00000000",
  1976 => x"00000000",
  1977 => x"00000000",
  1978 => x"00000000",
  1979 => x"25261e16",
  1980 => x"3e3d362e",
  1981 => x"48d0ff1e",
  1982 => x"7178e1c8",
  1983 => x"08d4ff48",
  1984 => x"1e4f2678",
  1985 => x"c848d0ff",
  1986 => x"487178e1",
  1987 => x"7808d4ff",
  1988 => x"ff4866c4",
  1989 => x"267808d4",
  1990 => x"4a711e4f",
  1991 => x"1e4966c4",
  1992 => x"deff4972",
  1993 => x"48d0ff87",
  1994 => x"2678e0c0",
  1995 => x"711e4f26",
  1996 => x"1e66c44a",
  1997 => x"49a2e0c1",
  1998 => x"c887c8ff",
  1999 => x"b7c84966",
  2000 => x"48d4ff29",
  2001 => x"d0ff7871",
  2002 => x"78e0c048",
  2003 => x"1e4f2626",
  2004 => x"c34ad4ff",
  2005 => x"d0ff7aff",
  2006 => x"78e1c848",
  2007 => x"cac47ade",
  2008 => x"497abff1",
  2009 => x"7028c848",
  2010 => x"d048717a",
  2011 => x"717a7028",
  2012 => x"7028d848",
  2013 => x"48d0ff7a",
  2014 => x"2678e0c0",
  2015 => x"5b5e0e4f",
  2016 => x"710e5d5c",
  2017 => x"f1cac44c",
  2018 => x"744b4dbf",
  2019 => x"9b66d02b",
  2020 => x"66d483c1",
  2021 => x"87c204ab",
  2022 => x"4a744bc0",
  2023 => x"724966d0",
  2024 => x"75b9ff31",
  2025 => x"72487399",
  2026 => x"484a7030",
  2027 => x"cac4b071",
  2028 => x"dafe58f5",
  2029 => x"264d2687",
  2030 => x"264b264c",
  2031 => x"d0ff1e4f",
  2032 => x"78c9c848",
  2033 => x"d4ff4871",
  2034 => x"4f267808",
  2035 => x"494a711e",
  2036 => x"d0ff87eb",
  2037 => x"2678c848",
  2038 => x"1e731e4f",
  2039 => x"cbc44b71",
  2040 => x"c302bfc1",
  2041 => x"87ebc287",
  2042 => x"c848d0ff",
  2043 => x"497378c9",
  2044 => x"ffb1e0c0",
  2045 => x"787148d4",
  2046 => x"48f5cac4",
  2047 => x"66c878c0",
  2048 => x"c387c502",
  2049 => x"87c249ff",
  2050 => x"cac449c0",
  2051 => x"66cc59fd",
  2052 => x"c587c602",
  2053 => x"c44ad5d5",
  2054 => x"ffffcf87",
  2055 => x"c1cbc44a",
  2056 => x"c1cbc45a",
  2057 => x"c478c148",
  2058 => x"264d2687",
  2059 => x"264b264c",
  2060 => x"5b5e0e4f",
  2061 => x"710e5d5c",
  2062 => x"fdcac44a",
  2063 => x"9a724cbf",
  2064 => x"4987cb02",
  2065 => x"ffc191c8",
  2066 => x"83714bcf",
  2067 => x"c3c287c4",
  2068 => x"4dc04bcf",
  2069 => x"99744913",
  2070 => x"bff9cac4",
  2071 => x"48d4ffb9",
  2072 => x"b7c17871",
  2073 => x"b7c8852c",
  2074 => x"87e804ad",
  2075 => x"bff5cac4",
  2076 => x"c480c848",
  2077 => x"fe58f9ca",
  2078 => x"731e87ef",
  2079 => x"134b711e",
  2080 => x"cb029a4a",
  2081 => x"fe497287",
  2082 => x"4a1387e7",
  2083 => x"87f5059a",
  2084 => x"1e87dafe",
  2085 => x"bff5cac4",
  2086 => x"f5cac449",
  2087 => x"78a1c148",
  2088 => x"a9b7c0c4",
  2089 => x"ff87db03",
  2090 => x"cac448d4",
  2091 => x"c478bff9",
  2092 => x"49bff5ca",
  2093 => x"48f5cac4",
  2094 => x"c478a1c1",
  2095 => x"04a9b7c0",
  2096 => x"d0ff87e5",
  2097 => x"c478c848",
  2098 => x"c048c1cb",
  2099 => x"004f2678",
  2100 => x"00000000",
  2101 => x"00000000",
  2102 => x"5f5f0000",
  2103 => x"00000000",
  2104 => x"03000303",
  2105 => x"14000003",
  2106 => x"7f147f7f",
  2107 => x"0000147f",
  2108 => x"6b6b2e24",
  2109 => x"4c00123a",
  2110 => x"6c18366a",
  2111 => x"30003256",
  2112 => x"77594f7e",
  2113 => x"0040683a",
  2114 => x"03070400",
  2115 => x"00000000",
  2116 => x"633e1c00",
  2117 => x"00000041",
  2118 => x"3e634100",
  2119 => x"0800001c",
  2120 => x"1c1c3e2a",
  2121 => x"00082a3e",
  2122 => x"3e3e0808",
  2123 => x"00000808",
  2124 => x"60e08000",
  2125 => x"00000000",
  2126 => x"08080808",
  2127 => x"00000808",
  2128 => x"60600000",
  2129 => x"40000000",
  2130 => x"0c183060",
  2131 => x"00010306",
  2132 => x"4d597f3e",
  2133 => x"00003e7f",
  2134 => x"7f7f0604",
  2135 => x"00000000",
  2136 => x"59716342",
  2137 => x"0000464f",
  2138 => x"49496322",
  2139 => x"1800367f",
  2140 => x"7f13161c",
  2141 => x"0000107f",
  2142 => x"45456727",
  2143 => x"0000397d",
  2144 => x"494b7e3c",
  2145 => x"00003079",
  2146 => x"79710101",
  2147 => x"0000070f",
  2148 => x"49497f36",
  2149 => x"0000367f",
  2150 => x"69494f06",
  2151 => x"00001e3f",
  2152 => x"66660000",
  2153 => x"00000000",
  2154 => x"66e68000",
  2155 => x"00000000",
  2156 => x"14140808",
  2157 => x"00002222",
  2158 => x"14141414",
  2159 => x"00001414",
  2160 => x"14142222",
  2161 => x"00000808",
  2162 => x"59510302",
  2163 => x"3e00060f",
  2164 => x"555d417f",
  2165 => x"00001e1f",
  2166 => x"09097f7e",
  2167 => x"00007e7f",
  2168 => x"49497f7f",
  2169 => x"0000367f",
  2170 => x"41633e1c",
  2171 => x"00004141",
  2172 => x"63417f7f",
  2173 => x"00001c3e",
  2174 => x"49497f7f",
  2175 => x"00004141",
  2176 => x"09097f7f",
  2177 => x"00000101",
  2178 => x"49417f3e",
  2179 => x"00007a7b",
  2180 => x"08087f7f",
  2181 => x"00007f7f",
  2182 => x"7f7f4100",
  2183 => x"00000041",
  2184 => x"40406020",
  2185 => x"7f003f7f",
  2186 => x"361c087f",
  2187 => x"00004163",
  2188 => x"40407f7f",
  2189 => x"7f004040",
  2190 => x"060c067f",
  2191 => x"7f007f7f",
  2192 => x"180c067f",
  2193 => x"00007f7f",
  2194 => x"41417f3e",
  2195 => x"00003e7f",
  2196 => x"09097f7f",
  2197 => x"3e00060f",
  2198 => x"7f61417f",
  2199 => x"0000407e",
  2200 => x"19097f7f",
  2201 => x"0000667f",
  2202 => x"594d6f26",
  2203 => x"0000327b",
  2204 => x"7f7f0101",
  2205 => x"00000101",
  2206 => x"40407f3f",
  2207 => x"00003f7f",
  2208 => x"70703f0f",
  2209 => x"7f000f3f",
  2210 => x"3018307f",
  2211 => x"41007f7f",
  2212 => x"1c1c3663",
  2213 => x"01416336",
  2214 => x"7c7c0603",
  2215 => x"61010306",
  2216 => x"474d5971",
  2217 => x"00004143",
  2218 => x"417f7f00",
  2219 => x"01000041",
  2220 => x"180c0603",
  2221 => x"00406030",
  2222 => x"7f414100",
  2223 => x"0800007f",
  2224 => x"0603060c",
  2225 => x"8000080c",
  2226 => x"80808080",
  2227 => x"00008080",
  2228 => x"07030000",
  2229 => x"00000004",
  2230 => x"54547420",
  2231 => x"0000787c",
  2232 => x"44447f7f",
  2233 => x"0000387c",
  2234 => x"44447c38",
  2235 => x"00000044",
  2236 => x"44447c38",
  2237 => x"00007f7f",
  2238 => x"54547c38",
  2239 => x"0000185c",
  2240 => x"057f7e04",
  2241 => x"00000005",
  2242 => x"a4a4bc18",
  2243 => x"00007cfc",
  2244 => x"04047f7f",
  2245 => x"0000787c",
  2246 => x"7d3d0000",
  2247 => x"00000040",
  2248 => x"fd808080",
  2249 => x"0000007d",
  2250 => x"38107f7f",
  2251 => x"0000446c",
  2252 => x"7f3f0000",
  2253 => x"7c000040",
  2254 => x"0c180c7c",
  2255 => x"0000787c",
  2256 => x"04047c7c",
  2257 => x"0000787c",
  2258 => x"44447c38",
  2259 => x"0000387c",
  2260 => x"2424fcfc",
  2261 => x"0000183c",
  2262 => x"24243c18",
  2263 => x"0000fcfc",
  2264 => x"04047c7c",
  2265 => x"0000080c",
  2266 => x"54545c48",
  2267 => x"00002074",
  2268 => x"447f3f04",
  2269 => x"00000044",
  2270 => x"40407c3c",
  2271 => x"00007c7c",
  2272 => x"60603c1c",
  2273 => x"3c001c3c",
  2274 => x"6030607c",
  2275 => x"44003c7c",
  2276 => x"3810386c",
  2277 => x"0000446c",
  2278 => x"60e0bc1c",
  2279 => x"00001c3c",
  2280 => x"5c746444",
  2281 => x"0000444c",
  2282 => x"773e0808",
  2283 => x"00004141",
  2284 => x"7f7f0000",
  2285 => x"00000000",
  2286 => x"3e774141",
  2287 => x"02000808",
  2288 => x"02030101",
  2289 => x"7f000102",
  2290 => x"7f7f7f7f",
  2291 => x"08007f7f",
  2292 => x"3e1c1c08",
  2293 => x"7f7f7f3e",
  2294 => x"1c3e3e7f",
  2295 => x"0008081c",
  2296 => x"7c7c1810",
  2297 => x"00001018",
  2298 => x"7c7c3010",
  2299 => x"10001030",
  2300 => x"78606030",
  2301 => x"4200061e",
  2302 => x"3c183c66",
  2303 => x"78004266",
  2304 => x"c6c26a38",
  2305 => x"6000386c",
  2306 => x"00600000",
  2307 => x"0e006000",
  2308 => x"5d5c5b5e",
  2309 => x"4c711e0e",
  2310 => x"bfd2cbc4",
  2311 => x"c04bc04d",
  2312 => x"02ab741e",
  2313 => x"a6c487c7",
  2314 => x"c578c048",
  2315 => x"48a6c487",
  2316 => x"66c478c1",
  2317 => x"ee49731e",
  2318 => x"86c887df",
  2319 => x"ef49e0c0",
  2320 => x"a5c487ef",
  2321 => x"f0496a4a",
  2322 => x"c6f187f0",
  2323 => x"c185cb87",
  2324 => x"abb7c883",
  2325 => x"87c7ff04",
  2326 => x"264d2626",
  2327 => x"264b264c",
  2328 => x"4a711e4f",
  2329 => x"5ad6cbc4",
  2330 => x"48d6cbc4",
  2331 => x"fe4978c7",
  2332 => x"4f2687dd",
  2333 => x"711e731e",
  2334 => x"aab7c04a",
  2335 => x"c287d303",
  2336 => x"05bfc8e0",
  2337 => x"4bc187c4",
  2338 => x"4bc087c2",
  2339 => x"5bcce0c2",
  2340 => x"e0c287c4",
  2341 => x"e0c25acc",
  2342 => x"c14abfc8",
  2343 => x"a2c0c19a",
  2344 => x"87e8ec49",
  2345 => x"e0c248fc",
  2346 => x"fe78bfc8",
  2347 => x"711e87ef",
  2348 => x"1e66c44a",
  2349 => x"f5e94972",
  2350 => x"4f262687",
  2351 => x"c8e0c21e",
  2352 => x"c8e649bf",
  2353 => x"cacbc487",
  2354 => x"78bfe848",
  2355 => x"48c6cbc4",
  2356 => x"c478bfec",
  2357 => x"4abfcacb",
  2358 => x"99ffcf49",
  2359 => x"722ab7ca",
  2360 => x"c4b07148",
  2361 => x"2658d2cb",
  2362 => x"5b5e0e4f",
  2363 => x"710e5d5c",
  2364 => x"87c8ff4b",
  2365 => x"48c5cbc4",
  2366 => x"497350c0",
  2367 => x"7087f5e5",
  2368 => x"9cc24c49",
  2369 => x"c149eecb",
  2370 => x"7087cfd7",
  2371 => x"cbc44d49",
  2372 => x"05bf97c5",
  2373 => x"d087e3c1",
  2374 => x"cbc44966",
  2375 => x"0599bfce",
  2376 => x"66d487d6",
  2377 => x"c6cbc449",
  2378 => x"cb0599bf",
  2379 => x"e5497387",
  2380 => x"987087c2",
  2381 => x"87c2c102",
  2382 => x"fffd4cc1",
  2383 => x"c1497587",
  2384 => x"7087e3d6",
  2385 => x"87c60298",
  2386 => x"48c5cbc4",
  2387 => x"cbc450c1",
  2388 => x"05bf97c5",
  2389 => x"c487e3c0",
  2390 => x"49bfcecb",
  2391 => x"059966d0",
  2392 => x"c487d5ff",
  2393 => x"49bfc6cb",
  2394 => x"059966d4",
  2395 => x"7387c9ff",
  2396 => x"87c0e449",
  2397 => x"fe059870",
  2398 => x"487487fe",
  2399 => x"0e87dafb",
  2400 => x"5d5c5b5e",
  2401 => x"c086f40e",
  2402 => x"bfec4c4d",
  2403 => x"48a6c47e",
  2404 => x"bfd2cbc4",
  2405 => x"c01ec178",
  2406 => x"fd49c71e",
  2407 => x"86c887cb",
  2408 => x"cd029870",
  2409 => x"fb49ff87",
  2410 => x"dac187ca",
  2411 => x"87c4e349",
  2412 => x"cbc44dc1",
  2413 => x"02bf97c5",
  2414 => x"e0c187c4",
  2415 => x"cbc487ff",
  2416 => x"c24bbfca",
  2417 => x"05bfc8e0",
  2418 => x"c487dac1",
  2419 => x"c0c248a6",
  2420 => x"c378c0c0",
  2421 => x"6e7ecff9",
  2422 => x"6e49bf97",
  2423 => x"7080c148",
  2424 => x"cfe2717e",
  2425 => x"02987087",
  2426 => x"66c487c3",
  2427 => x"4866c4b3",
  2428 => x"c828b7c1",
  2429 => x"987058a6",
  2430 => x"87dbff05",
  2431 => x"e149fdc3",
  2432 => x"fac387f2",
  2433 => x"87ece149",
  2434 => x"ffcf4973",
  2435 => x"c01e7199",
  2436 => x"87dafa49",
  2437 => x"b7ca4973",
  2438 => x"c11e7129",
  2439 => x"87cefa49",
  2440 => x"c7c686c8",
  2441 => x"cecbc487",
  2442 => x"029b4bbf",
  2443 => x"e0c287df",
  2444 => x"c149bfc4",
  2445 => x"7087efd2",
  2446 => x"87c40598",
  2447 => x"87d34bc0",
  2448 => x"c149e0c2",
  2449 => x"c287d3d2",
  2450 => x"c658c8e0",
  2451 => x"c4e0c287",
  2452 => x"7378c048",
  2453 => x"0599c249",
  2454 => x"ebc387ce",
  2455 => x"87d4e049",
  2456 => x"99c24970",
  2457 => x"87c2c002",
  2458 => x"49734cfb",
  2459 => x"cf0599c1",
  2460 => x"49f4c387",
  2461 => x"87fcdfff",
  2462 => x"99c24970",
  2463 => x"87c2c002",
  2464 => x"49734cfa",
  2465 => x"ce0599c8",
  2466 => x"49f5c387",
  2467 => x"87e4dfff",
  2468 => x"99c24970",
  2469 => x"c487d602",
  2470 => x"02bfd6cb",
  2471 => x"4887cac0",
  2472 => x"cbc488c1",
  2473 => x"c2c058da",
  2474 => x"c14cff87",
  2475 => x"c449734d",
  2476 => x"cec00599",
  2477 => x"49f2c387",
  2478 => x"87f8deff",
  2479 => x"99c24970",
  2480 => x"c487dc02",
  2481 => x"7ebfd6cb",
  2482 => x"a8b7c748",
  2483 => x"87cbc003",
  2484 => x"80c1486e",
  2485 => x"58dacbc4",
  2486 => x"fe87c2c0",
  2487 => x"c34dc14c",
  2488 => x"deff49fd",
  2489 => x"497087ce",
  2490 => x"c00299c2",
  2491 => x"cbc487d5",
  2492 => x"c002bfd6",
  2493 => x"cbc487c9",
  2494 => x"78c048d6",
  2495 => x"fd87c2c0",
  2496 => x"c34dc14c",
  2497 => x"ddff49fa",
  2498 => x"497087ea",
  2499 => x"c00299c2",
  2500 => x"cbc487d9",
  2501 => x"c748bfd6",
  2502 => x"c003a8b7",
  2503 => x"cbc487c9",
  2504 => x"78c748d6",
  2505 => x"fc87c2c0",
  2506 => x"c04dc14c",
  2507 => x"c003acb7",
  2508 => x"66c487d1",
  2509 => x"82d8c14a",
  2510 => x"c6c0026a",
  2511 => x"744b6a87",
  2512 => x"c00f7349",
  2513 => x"1ef0c31e",
  2514 => x"f649dac1",
  2515 => x"86c887db",
  2516 => x"c0029870",
  2517 => x"a6c887e2",
  2518 => x"d6cbc448",
  2519 => x"66c878bf",
  2520 => x"c491cb49",
  2521 => x"80714866",
  2522 => x"bf6e7e70",
  2523 => x"87c8c002",
  2524 => x"c84bbf6e",
  2525 => x"0f734966",
  2526 => x"c0029d75",
  2527 => x"cbc487c8",
  2528 => x"f249bfd6",
  2529 => x"e0c287c9",
  2530 => x"c002bfcc",
  2531 => x"c14987de",
  2532 => x"7087d3cd",
  2533 => x"d3c00298",
  2534 => x"d6cbc487",
  2535 => x"eef149bf",
  2536 => x"f349c087",
  2537 => x"e0c287ce",
  2538 => x"78c048cc",
  2539 => x"e8f28ef4",
  2540 => x"5b5e0e87",
  2541 => x"1e0e5d5c",
  2542 => x"cbc44c71",
  2543 => x"c149bfd2",
  2544 => x"c14da1cd",
  2545 => x"7e6981d1",
  2546 => x"cf029c74",
  2547 => x"4ba5c487",
  2548 => x"cbc47b74",
  2549 => x"f249bfd2",
  2550 => x"7b6e87c7",
  2551 => x"c4059c74",
  2552 => x"c24bc087",
  2553 => x"734bc187",
  2554 => x"87c8f249",
  2555 => x"c90266d4",
  2556 => x"cbc14987",
  2557 => x"4a7087e4",
  2558 => x"4ac087c2",
  2559 => x"5ad0e0c2",
  2560 => x"87d5f126",
  2561 => x"00000000",
  2562 => x"00000000",
  2563 => x"00000000",
  2564 => x"711e731e",
  2565 => x"cbc1494b",
  2566 => x"f6e8fd4a",
  2567 => x"1e4a7087",
  2568 => x"fcc04972",
  2569 => x"eae8fd4a",
  2570 => x"26497087",
  2571 => x"4866c84a",
  2572 => x"49725071",
  2573 => x"fd4afcc0",
  2574 => x"7187d8e8",
  2575 => x"4966c84a",
  2576 => x"517281c1",
  2577 => x"cbc14973",
  2578 => x"c6e8fd4a",
  2579 => x"c84a7187",
  2580 => x"81c24966",
  2581 => x"87c45172",
  2582 => x"4c264d26",
  2583 => x"4f264b26",
  2584 => x"711e731e",
  2585 => x"4966c84b",
  2586 => x"cc91cbc1",
  2587 => x"49a14a66",
  2588 => x"c6c14a73",
  2589 => x"a17292d4",
  2590 => x"89d6c249",
  2591 => x"dbff4871",
  2592 => x"5b5e0e87",
  2593 => x"1e0e5d5c",
  2594 => x"6b974b71",
  2595 => x"87e4c002",
  2596 => x"487e6b97",
  2597 => x"a8b7f0c0",
  2598 => x"6e87d904",
  2599 => x"b7f9c048",
  2600 => x"87d001a8",
  2601 => x"496e83c1",
  2602 => x"ca89f0c0",
  2603 => x"4866d491",
  2604 => x"87c55071",
  2605 => x"ebc448c0",
  2606 => x"026b9787",
  2607 => x"9787e9c0",
  2608 => x"c0487e6b",
  2609 => x"04a8b7f0",
  2610 => x"486e87de",
  2611 => x"a8b7f9c0",
  2612 => x"c187d501",
  2613 => x"c0496e83",
  2614 => x"66d489f0",
  2615 => x"a14abf97",
  2616 => x"4866d449",
  2617 => x"87c55071",
  2618 => x"f7c348c0",
  2619 => x"026b9787",
  2620 => x"6b9787cd",
  2621 => x"a9fac049",
  2622 => x"c187c405",
  2623 => x"c087c583",
  2624 => x"87e0c348",
  2625 => x"c0026b97",
  2626 => x"6b9787e7",
  2627 => x"f0c0487e",
  2628 => x"dc04a8b7",
  2629 => x"c0486e87",
  2630 => x"01a8b7f9",
  2631 => x"83c187d3",
  2632 => x"f0c0496e",
  2633 => x"d491ca89",
  2634 => x"84c14c66",
  2635 => x"c57c9771",
  2636 => x"c248c087",
  2637 => x"6b9787ee",
  2638 => x"87e4c002",
  2639 => x"487e6b97",
  2640 => x"a8b7f0c0",
  2641 => x"6e87d904",
  2642 => x"b7f9c048",
  2643 => x"87d001a8",
  2644 => x"496e83c1",
  2645 => x"9789f0c0",
  2646 => x"49a14a6c",
  2647 => x"87c57c97",
  2648 => x"ffc148c0",
  2649 => x"026b9787",
  2650 => x"6b9787cd",
  2651 => x"a9fac049",
  2652 => x"c187c405",
  2653 => x"c087c583",
  2654 => x"87e8c148",
  2655 => x"c0026b97",
  2656 => x"6b9787e4",
  2657 => x"b7f0c04a",
  2658 => x"87da04aa",
  2659 => x"aab7f9c0",
  2660 => x"c187d301",
  2661 => x"c0497283",
  2662 => x"91ca89f0",
  2663 => x"c24d66d4",
  2664 => x"7d977185",
  2665 => x"48c087c5",
  2666 => x"9787f9c0",
  2667 => x"e4c0026b",
  2668 => x"7e6b9787",
  2669 => x"b7f0c048",
  2670 => x"87d904a8",
  2671 => x"f9c0486e",
  2672 => x"d001a8b7",
  2673 => x"6e83c187",
  2674 => x"89f0c049",
  2675 => x"a14a6d97",
  2676 => x"c47d9749",
  2677 => x"cb48c087",
  2678 => x"026b9787",
  2679 => x"48c087c4",
  2680 => x"48c187c2",
  2681 => x"87f0f926",
  2682 => x"5c5b5e0e",
  2683 => x"86f80e5d",
  2684 => x"4cc04d71",
  2685 => x"d2ccc44b",
  2686 => x"eecbfe49",
  2687 => x"c04a7087",
  2688 => x"c204aab7",
  2689 => x"aaca87f2",
  2690 => x"87ecc202",
  2691 => x"02aae0c0",
  2692 => x"aac987cf",
  2693 => x"cd87ca02",
  2694 => x"87c502aa",
  2695 => x"c605aaca",
  2696 => x"029c7487",
  2697 => x"c087d1c2",
  2698 => x"cc05aae2",
  2699 => x"c1497487",
  2700 => x"c34c71b9",
  2701 => x"fcfe9cff",
  2702 => x"059c7487",
  2703 => x"c187e7c1",
  2704 => x"04aab7e1",
  2705 => x"fac187c8",
  2706 => x"c106aab7",
  2707 => x"c1c187d8",
  2708 => x"c804aab7",
  2709 => x"b7dac187",
  2710 => x"c9c106aa",
  2711 => x"b7f0c087",
  2712 => x"87c804aa",
  2713 => x"aab7f9c0",
  2714 => x"87fac006",
  2715 => x"02aadbc1",
  2716 => x"c187f3c0",
  2717 => x"c002aadd",
  2718 => x"edc087ec",
  2719 => x"e5c002aa",
  2720 => x"aadfc187",
  2721 => x"c087df02",
  2722 => x"d902aaec",
  2723 => x"aafdc087",
  2724 => x"c187d302",
  2725 => x"cd02aafe",
  2726 => x"aafac087",
  2727 => x"c087c702",
  2728 => x"fd05aaef",
  2729 => x"ffc087cf",
  2730 => x"fd03abb7",
  2731 => x"a37587c7",
  2732 => x"7283c149",
  2733 => x"87fdfc51",
  2734 => x"c049a375",
  2735 => x"03aab751",
  2736 => x"7ec487c4",
  2737 => x"9b7387df",
  2738 => x"c487c705",
  2739 => x"78c348a6",
  2740 => x"9c7487d0",
  2741 => x"c187c402",
  2742 => x"c087c27e",
  2743 => x"48a6c47e",
  2744 => x"66c4786e",
  2745 => x"f8486e7e",
  2746 => x"87ecf58e",
  2747 => x"5c5b5e0e",
  2748 => x"4d710e5d",
  2749 => x"4bdacbc4",
  2750 => x"f8c04ac0",
  2751 => x"d5d7fd49",
  2752 => x"c41e7587",
  2753 => x"fd49d2cc",
  2754 => x"c487c3fc",
  2755 => x"05987086",
  2756 => x"4cc187c5",
  2757 => x"c187eac0",
  2758 => x"87eac049",
  2759 => x"059c4c70",
  2760 => x"cbc487c9",
  2761 => x"dd49bfde",
  2762 => x"744c7087",
  2763 => x"87cb059c",
  2764 => x"48dacbc4",
  2765 => x"bfeecbc4",
  2766 => x"c487c678",
  2767 => x"c048decb",
  2768 => x"f4487478",
  2769 => x"5e0e87d2",
  2770 => x"0e5d5c5b",
  2771 => x"7186d4ff",
  2772 => x"7e97c04c",
  2773 => x"c048a6c4",
  2774 => x"5080c050",
  2775 => x"c05080c0",
  2776 => x"c04d5080",
  2777 => x"80c47880",
  2778 => x"80c478c0",
  2779 => x"80c478c0",
  2780 => x"ccc478c0",
  2781 => x"c505bfda",
  2782 => x"d048c187",
  2783 => x"ccc487c3",
  2784 => x"78c048d2",
  2785 => x"78c080d0",
  2786 => x"ccc480f4",
  2787 => x"c378bfde",
  2788 => x"c048f3c0",
  2789 => x"eecbc478",
  2790 => x"c278c048",
  2791 => x"f949f3ff",
  2792 => x"a6dc87c6",
  2793 => x"02a8c358",
  2794 => x"9787d0cd",
  2795 => x"029b4b6e",
  2796 => x"8bc187d8",
  2797 => x"87f5c102",
  2798 => x"e4c3028b",
  2799 => x"c7028b87",
  2800 => x"028b87c4",
  2801 => x"cc87c3c8",
  2802 => x"a6c487f1",
  2803 => x"c250c048",
  2804 => x"c24af3ff",
  2805 => x"fd49e3fe",
  2806 => x"7087f4d1",
  2807 => x"87c60598",
  2808 => x"cc7e97c1",
  2809 => x"ffc287d5",
  2810 => x"fec24af3",
  2811 => x"d1fd49e8",
  2812 => x"987087dd",
  2813 => x"c287c605",
  2814 => x"fecb7e97",
  2815 => x"f3ffc287",
  2816 => x"eefec24a",
  2817 => x"c6d1fd49",
  2818 => x"05987087",
  2819 => x"c387c6c0",
  2820 => x"e6cb7e97",
  2821 => x"f3ffc287",
  2822 => x"f5fec24a",
  2823 => x"eed0fd49",
  2824 => x"05987087",
  2825 => x"c487d4cb",
  2826 => x"cecb7e97",
  2827 => x"6697c487",
  2828 => x"a6e0c048",
  2829 => x"05987058",
  2830 => x"c887cdc1",
  2831 => x"78c048a6",
  2832 => x"056697c7",
  2833 => x"c487cdc1",
  2834 => x"02bfc6cc",
  2835 => x"ff87c7c0",
  2836 => x"c050c180",
  2837 => x"ffc287fe",
  2838 => x"cbc41ef3",
  2839 => x"f6fd49fe",
  2840 => x"86c487ec",
  2841 => x"c0029870",
  2842 => x"a6c787c8",
  2843 => x"c050c148",
  2844 => x"a6c587c5",
  2845 => x"c350c448",
  2846 => x"c41ecafa",
  2847 => x"fd49d2cc",
  2848 => x"c487e7f9",
  2849 => x"87ccc086",
  2850 => x"c14866dc",
  2851 => x"c3c005a8",
  2852 => x"7e97c087",
  2853 => x"486697c4",
  2854 => x"a6c480c1",
  2855 => x"dac95008",
  2856 => x"48a6d487",
  2857 => x"7866e0c0",
  2858 => x"486697c4",
  2859 => x"58a6e0c0",
  2860 => x"c0059870",
  2861 => x"1eca87fb",
  2862 => x"ffc21ec0",
  2863 => x"d3fd49f3",
  2864 => x"86c887cf",
  2865 => x"e0c04970",
  2866 => x"66dc59a6",
  2867 => x"87d3c002",
  2868 => x"b7e3c148",
  2869 => x"cac001a8",
  2870 => x"49a5c187",
  2871 => x"02a966dc",
  2872 => x"c587c8c0",
  2873 => x"50c248a6",
  2874 => x"dc87cec2",
  2875 => x"c8c24d66",
  2876 => x"4866dc87",
  2877 => x"c105a8c1",
  2878 => x"ffc287ff",
  2879 => x"fec24af3",
  2880 => x"cdfd49c7",
  2881 => x"987087c9",
  2882 => x"87cfc005",
  2883 => x"48a6e0c0",
  2884 => x"78f0e4c0",
  2885 => x"78c080c4",
  2886 => x"c287c7c1",
  2887 => x"c24af3ff",
  2888 => x"fd49cdfe",
  2889 => x"7087e8cc",
  2890 => x"cfc00598",
  2891 => x"a6e0c087",
  2892 => x"f0e4c048",
  2893 => x"c180c478",
  2894 => x"87e6c078",
  2895 => x"4af3ffc2",
  2896 => x"49d8fec2",
  2897 => x"87c7ccfd",
  2898 => x"c0059870",
  2899 => x"e0c087cf",
  2900 => x"e0c048a6",
  2901 => x"80c478c0",
  2902 => x"c5c078c1",
  2903 => x"48a6c587",
  2904 => x"ac7550c2",
  2905 => x"87cec005",
  2906 => x"48f6cbc4",
  2907 => x"7866e0c0",
  2908 => x"e4c080fc",
  2909 => x"97c07866",
  2910 => x"6697c47e",
  2911 => x"c480c148",
  2912 => x"c55008a6",
  2913 => x"e8c087f5",
  2914 => x"ffc21ea6",
  2915 => x"f0eb49f3",
  2916 => x"7086c487",
  2917 => x"c8c00598",
  2918 => x"48a6c587",
  2919 => x"e3c050c2",
  2920 => x"97eac087",
  2921 => x"c01e4966",
  2922 => x"496697ed",
  2923 => x"97f0c01e",
  2924 => x"ebea4966",
  2925 => x"7086c887",
  2926 => x"81d6c249",
  2927 => x"66c84871",
  2928 => x"58a6cc80",
  2929 => x"c47e97c0",
  2930 => x"97c487f1",
  2931 => x"e0c04866",
  2932 => x"987058a6",
  2933 => x"87d7c005",
  2934 => x"1ec01eca",
  2935 => x"49f3ffc2",
  2936 => x"87edcefd",
  2937 => x"497086c8",
  2938 => x"5997a6ca",
  2939 => x"dc87c2c4",
  2940 => x"a8c14866",
  2941 => x"87f9c305",
  2942 => x"1ea6e8c0",
  2943 => x"49f3ffc2",
  2944 => x"c487fee9",
  2945 => x"05987086",
  2946 => x"c587c8c0",
  2947 => x"50c248a6",
  2948 => x"c087dbc3",
  2949 => x"496697ea",
  2950 => x"97edc01e",
  2951 => x"c01e4966",
  2952 => x"496697f0",
  2953 => x"c887f9e8",
  2954 => x"c67e7086",
  2955 => x"c0486697",
  2956 => x"7058a6e0",
  2957 => x"e1c00598",
  2958 => x"49a4c187",
  2959 => x"edc205ad",
  2960 => x"eecbc487",
  2961 => x"e5c205bf",
  2962 => x"c2496e87",
  2963 => x"487181d6",
  2964 => x"c48066c8",
  2965 => x"c258f2cb",
  2966 => x"66dc87d4",
  2967 => x"05a8c148",
  2968 => x"7487cbc2",
  2969 => x"cec005ad",
  2970 => x"c2496e87",
  2971 => x"487181d6",
  2972 => x"c48066c8",
  2973 => x"c158eecb",
  2974 => x"c106adb7",
  2975 => x"486e87ce",
  2976 => x"c08866cc",
  2977 => x"7458a6e0",
  2978 => x"cec005ad",
  2979 => x"d4497087",
  2980 => x"48719166",
  2981 => x"c48066d0",
  2982 => x"c158eacb",
  2983 => x"05ad49a4",
  2984 => x"c487d8c0",
  2985 => x"05bfeecb",
  2986 => x"6e87d0c0",
  2987 => x"81d6c249",
  2988 => x"718166c8",
  2989 => x"c488c148",
  2990 => x"dc58f2cb",
  2991 => x"66d44966",
  2992 => x"d0487191",
  2993 => x"a6d48066",
  2994 => x"87ddc058",
  2995 => x"d6c2496e",
  2996 => x"9166d481",
  2997 => x"66d04871",
  2998 => x"58a6d480",
  2999 => x"c005acc1",
  3000 => x"cbc487c7",
  3001 => x"66d048e6",
  3002 => x"48a6cc78",
  3003 => x"97c0786e",
  3004 => x"6697c47e",
  3005 => x"c480c148",
  3006 => x"d85008a6",
  3007 => x"a8c44866",
  3008 => x"87c7c002",
  3009 => x"026697c5",
  3010 => x"c787d0f2",
  3011 => x"c0056697",
  3012 => x"a6c587c8",
  3013 => x"c050c448",
  3014 => x"ad7487f1",
  3015 => x"87ebc005",
  3016 => x"bfe6cbc4",
  3017 => x"c6ccc44a",
  3018 => x"887248bf",
  3019 => x"cbc44a70",
  3020 => x"7249bff6",
  3021 => x"4a09721e",
  3022 => x"87e3cbfd",
  3023 => x"4a264970",
  3024 => x"bfeacbc4",
  3025 => x"c4807148",
  3026 => x"7458f2cb",
  3027 => x"c003adb7",
  3028 => x"a6c587c5",
  3029 => x"c550c448",
  3030 => x"c0026697",
  3031 => x"cbc487c9",
  3032 => x"78c048de",
  3033 => x"c487c4c0",
  3034 => x"c05de2cb",
  3035 => x"c41ea6e8",
  3036 => x"49bfeacb",
  3037 => x"c487d9e2",
  3038 => x"fecbc486",
  3039 => x"6697c55c",
  3040 => x"8ed4ff48",
  3041 => x"4187d1e3",
  3042 => x"4f494455",
  3043 => x"444f4d00",
  3044 => x"322f3145",
  3045 => x"00323533",
  3046 => x"45444f4d",
  3047 => x"30322f31",
  3048 => x"46003834",
  3049 => x"00454c49",
  3050 => x"43415254",
  3051 => x"5250004b",
  3052 => x"50414745",
  3053 => x"444e4900",
  3054 => x"0e005845",
  3055 => x"0e5c5b5e",
  3056 => x"4cc14b71",
  3057 => x"bfeacbc4",
  3058 => x"d004abb7",
  3059 => x"eecbc487",
  3060 => x"01abb7bf",
  3061 => x"cbc487c7",
  3062 => x"d348bffa",
  3063 => x"ed497487",
  3064 => x"84c187e4",
  3065 => x"bfdecbc4",
  3066 => x"ff06acb7",
  3067 => x"48ff87d6",
  3068 => x"0087e7e1",
  3069 => x"00000000",
  3070 => x"00000000",
  3071 => x"00000000",
  3072 => x"00000000",
  3073 => x"00000000",
  3074 => x"00000000",
  3075 => x"00000000",
  3076 => x"00000000",
  3077 => x"00000000",
  3078 => x"00000000",
  3079 => x"00000000",
  3080 => x"00000000",
  3081 => x"00000000",
  3082 => x"00000000",
  3083 => x"00000000",
  3084 => x"00000000",
  3085 => x"1e000000",
  3086 => x"4b711e73",
  3087 => x"49721e4a",
  3088 => x"c8fd4aca",
  3089 => x"497087cd",
  3090 => x"91d04a26",
  3091 => x"49721e71",
  3092 => x"c7fd4aca",
  3093 => x"4a7187fd",
  3094 => x"a1724926",
  3095 => x"99ffc349",
  3096 => x"87c44871",
  3097 => x"4c264d26",
  3098 => x"4f264b26",
  3099 => x"711e731e",
  3100 => x"c4494a4b",
  3101 => x"91ca29b7",
  3102 => x"a1729acf",
  3103 => x"99ffc349",
  3104 => x"87e44871",
  3105 => x"711e731e",
  3106 => x"87e0494a",
  3107 => x"9b4b4970",
  3108 => x"c187c205",
  3109 => x"decbc44b",
  3110 => x"06abb7bf",
  3111 => x"734b87c1",
  3112 => x"87e2ea49",
  3113 => x"fffe4873",
  3114 => x"f1c41e87",
  3115 => x"c45997da",
  3116 => x"c448d7f1",
  3117 => x"66c85066",
  3118 => x"5066cc50",
  3119 => x"731e4f26",
  3120 => x"ff4b711e",
  3121 => x"c5c848d0",
  3122 => x"48d4ff78",
  3123 => x"7378e1c1",
  3124 => x"b7c84a49",
  3125 => x"c378722a",
  3126 => x"787199ff",
  3127 => x"c448d0ff",
  3128 => x"87c4fe78",
  3129 => x"d4f2c41e",
  3130 => x"f1c4599f",
  3131 => x"78c148e4",
  3132 => x"5e0e4f26",
  3133 => x"710e5c5b",
  3134 => x"48d0ff4c",
  3135 => x"ff78c5c8",
  3136 => x"e4c148d4",
  3137 => x"4966cc78",
  3138 => x"9affc34a",
  3139 => x"66cc7872",
  3140 => x"c32ac84a",
  3141 => x"66d09aff",
  3142 => x"7333c74b",
  3143 => x"717872b2",
  3144 => x"fd49741e",
  3145 => x"ff87ddc5",
  3146 => x"78c448d0",
  3147 => x"87f6fc26",
  3148 => x"c01e731e",
  3149 => x"c44bc0e0",
  3150 => x"02bff2cb",
  3151 => x"c487e7c1",
  3152 => x"48bfeff1",
  3153 => x"04a8b7c0",
  3154 => x"c487dbc1",
  3155 => x"abbff6cb",
  3156 => x"c487d302",
  3157 => x"49bfcecc",
  3158 => x"1e7181d0",
  3159 => x"49fecbc4",
  3160 => x"87cce8fd",
  3161 => x"1e7386c4",
  3162 => x"1ee6ccc4",
  3163 => x"49fecbc4",
  3164 => x"87e3e9fd",
  3165 => x"cbc486c8",
  3166 => x"02abbff6",
  3167 => x"c04987d6",
  3168 => x"c489d0e0",
  3169 => x"81bfcecc",
  3170 => x"cbc41e71",
  3171 => x"e7fd49fe",
  3172 => x"86c487de",
  3173 => x"1e4966c8",
  3174 => x"ccc41e73",
  3175 => x"d1fd49e6",
  3176 => x"c086c887",
  3177 => x"e4c087e1",
  3178 => x"ccc41ef0",
  3179 => x"cbc41ee6",
  3180 => x"e8fd49fe",
  3181 => x"66d087e1",
  3182 => x"e4c01e49",
  3183 => x"ccc41ef0",
  3184 => x"edfc49e6",
  3185 => x"fa86d087",
  3186 => x"c41e87de",
  3187 => x"05bfc6cc",
  3188 => x"f1c487db",
  3189 => x"50c148de",
  3190 => x"cb1e1ec0",
  3191 => x"fb49c21e",
  3192 => x"86cc87c7",
  3193 => x"d5fb49c1",
  3194 => x"c248c087",
  3195 => x"2648c187",
  3196 => x"1e731e4f",
  3197 => x"bfdaf1c4",
  3198 => x"06a8c048",
  3199 => x"c387e9c0",
  3200 => x"49bfd6eb",
  3201 => x"87dee3c0",
  3202 => x"c7029870",
  3203 => x"49cd87e3",
  3204 => x"87c6e3c0",
  3205 => x"ebc34970",
  3206 => x"f1c459da",
  3207 => x"c148bfda",
  3208 => x"def1c488",
  3209 => x"87c9c758",
  3210 => x"97def1c4",
  3211 => x"aac24abf",
  3212 => x"87cac305",
  3213 => x"bfebf1c4",
  3214 => x"decbc448",
  3215 => x"06a8b7bf",
  3216 => x"f1c487c9",
  3217 => x"50c048de",
  3218 => x"c487e6c6",
  3219 => x"bf97e9f1",
  3220 => x"87ddc602",
  3221 => x"bfc6ccc4",
  3222 => x"c487da05",
  3223 => x"c148def1",
  3224 => x"1e1ec050",
  3225 => x"49c21ecb",
  3226 => x"cc87fef8",
  3227 => x"f949c186",
  3228 => x"fcc587f2",
  3229 => x"e9f1c487",
  3230 => x"c450c048",
  3231 => x"02bff2cb",
  3232 => x"1ec187cd",
  3233 => x"49c0e0c0",
  3234 => x"c487e5fa",
  3235 => x"c487d586",
  3236 => x"48bfeff1",
  3237 => x"bfeacbc4",
  3238 => x"c004a8b7",
  3239 => x"f1c487c6",
  3240 => x"50c048df",
  3241 => x"bff3f1c4",
  3242 => x"c488c148",
  3243 => x"7058f7f1",
  3244 => x"cbc00598",
  3245 => x"f849c087",
  3246 => x"f1c487ea",
  3247 => x"50c048de",
  3248 => x"bfeff1c4",
  3249 => x"c480c148",
  3250 => x"c458f3f1",
  3251 => x"b7bfeecb",
  3252 => x"dcc404a8",
  3253 => x"ebf1c487",
  3254 => x"80c148bf",
  3255 => x"58eff1c4",
  3256 => x"e1e14970",
  3257 => x"dff1c487",
  3258 => x"c450c148",
  3259 => x"49bfe6cb",
  3260 => x"fecbc41e",
  3261 => x"f7e1fd49",
  3262 => x"c386c487",
  3263 => x"aac387f3",
  3264 => x"87edc305",
  3265 => x"bfc6ccc4",
  3266 => x"87dac005",
  3267 => x"48def1c4",
  3268 => x"1ec050c1",
  3269 => x"c21ecb1e",
  3270 => x"87cdf649",
  3271 => x"49c186cc",
  3272 => x"c387c1f7",
  3273 => x"f1c487cb",
  3274 => x"f249bfef",
  3275 => x"f1c487cd",
  3276 => x"f1c458ef",
  3277 => x"05bf97ea",
  3278 => x"c087d5c1",
  3279 => x"cbf2c44b",
  3280 => x"b7c048bf",
  3281 => x"c7c104a8",
  3282 => x"f2cbc487",
  3283 => x"e8c005bf",
  3284 => x"eff1c487",
  3285 => x"cbc449bf",
  3286 => x"c089bfea",
  3287 => x"c491f0e4",
  3288 => x"81bfe6cb",
  3289 => x"cbc41e71",
  3290 => x"e0fd49fe",
  3291 => x"1ec087c2",
  3292 => x"49f0e4c0",
  3293 => x"c887f9f6",
  3294 => x"eff1c486",
  3295 => x"80c148bf",
  3296 => x"58f3f1c4",
  3297 => x"f2c483c1",
  3298 => x"abb7bfcb",
  3299 => x"87f9fe06",
  3300 => x"48cbf2c4",
  3301 => x"f1c478c0",
  3302 => x"c448bfef",
  3303 => x"b7bfc7f2",
  3304 => x"d7c003a8",
  3305 => x"f2cbc487",
  3306 => x"cfc005bf",
  3307 => x"ebf1c487",
  3308 => x"cbc448bf",
  3309 => x"a8b7bfde",
  3310 => x"87f5c006",
  3311 => x"97cff2c4",
  3312 => x"a9c149bf",
  3313 => x"87d2c005",
  3314 => x"48eff1c4",
  3315 => x"bfc3f2c4",
  3316 => x"daf1c478",
  3317 => x"c078c248",
  3318 => x"f1c487c6",
  3319 => x"50c048de",
  3320 => x"97cff2c4",
  3321 => x"a9c249bf",
  3322 => x"87c5c005",
  3323 => x"f3f349c0",
  3324 => x"87f4f187",
  3325 => x"5c5b5e0e",
  3326 => x"c4ff0e5d",
  3327 => x"c04b7686",
  3328 => x"49e0c04a",
  3329 => x"87cef3fc",
  3330 => x"c848d0ff",
  3331 => x"d4ff78c5",
  3332 => x"78e2c148",
  3333 => x"48a6e0c0",
  3334 => x"d4ff78c0",
  3335 => x"c078c048",
  3336 => x"c049a6e4",
  3337 => x"688166e0",
  3338 => x"66e0c051",
  3339 => x"c080c148",
  3340 => x"cc58a6e4",
  3341 => x"ff04a8b7",
  3342 => x"d0ff87e0",
  3343 => x"c078c448",
  3344 => x"4c6697e4",
  3345 => x"f3c0029c",
  3346 => x"028cc387",
  3347 => x"c587fec0",
  3348 => x"e5c6028c",
  3349 => x"028ccd87",
  3350 => x"c387e9c8",
  3351 => x"c8028cc3",
  3352 => x"8cc187fb",
  3353 => x"87d2cc02",
  3354 => x"c9d0028c",
  3355 => x"028cc387",
  3356 => x"c187dad0",
  3357 => x"f8c1028c",
  3358 => x"87ccd487",
  3359 => x"7087cbf5",
  3360 => x"ddd40298",
  3361 => x"f049c087",
  3362 => x"d5d487f4",
  3363 => x"7e97d287",
  3364 => x"c248a6c1",
  3365 => x"f0c150c0",
  3366 => x"c480c150",
  3367 => x"bf97d6f1",
  3368 => x"ca80c450",
  3369 => x"c480c450",
  3370 => x"bf97d7f1",
  3371 => x"d8f1c450",
  3372 => x"c450bf97",
  3373 => x"bf97d9f1",
  3374 => x"d9f1c450",
  3375 => x"c450c048",
  3376 => x"c448d8f1",
  3377 => x"bf97d9f1",
  3378 => x"d7f1c450",
  3379 => x"d8f1c448",
  3380 => x"c450bf97",
  3381 => x"c448d6f1",
  3382 => x"bf97d7f1",
  3383 => x"d21ec150",
  3384 => x"49a6ca1e",
  3385 => x"c887cbf0",
  3386 => x"ef49c086",
  3387 => x"f1d287d0",
  3388 => x"87d6f387",
  3389 => x"d2029870",
  3390 => x"e5c087e8",
  3391 => x"c0486697",
  3392 => x"7058a6e4",
  3393 => x"87da0298",
  3394 => x"c088c148",
  3395 => x"7058a6e4",
  3396 => x"edc00298",
  3397 => x"88c14887",
  3398 => x"58a6e4c0",
  3399 => x"c1029870",
  3400 => x"97c287eb",
  3401 => x"48a6c17e",
  3402 => x"c150c0c2",
  3403 => x"decbc450",
  3404 => x"c2ec49bf",
  3405 => x"08a6c387",
  3406 => x"a6e0c050",
  3407 => x"c278c248",
  3408 => x"cbc487e2",
  3409 => x"c249bfda",
  3410 => x"f0c081d6",
  3411 => x"ff711ea6",
  3412 => x"c487fdca",
  3413 => x"c17e9786",
  3414 => x"c0c248a6",
  3415 => x"97f0c050",
  3416 => x"d2eb4966",
  3417 => x"08a6c287",
  3418 => x"97f1c050",
  3419 => x"c6eb4966",
  3420 => x"08a6c387",
  3421 => x"97f2c050",
  3422 => x"faea4966",
  3423 => x"08a6c487",
  3424 => x"48a6c550",
  3425 => x"80da50c0",
  3426 => x"d7c178c4",
  3427 => x"97e6c087",
  3428 => x"efeb4966",
  3429 => x"eacbc487",
  3430 => x"d6c249bf",
  3431 => x"a6f0c081",
  3432 => x"c9ff711e",
  3433 => x"86c487ea",
  3434 => x"a6c17e97",
  3435 => x"50c0c248",
  3436 => x"6697f0c0",
  3437 => x"87ffe949",
  3438 => x"5008a6c2",
  3439 => x"6697f1c0",
  3440 => x"87f3e949",
  3441 => x"5008a6c3",
  3442 => x"6697f2c0",
  3443 => x"87e7e949",
  3444 => x"5008a6c4",
  3445 => x"bff2cbc4",
  3446 => x"c931c249",
  3447 => x"485997a6",
  3448 => x"78c480db",
  3449 => x"e4c01ec1",
  3450 => x"a6ca1e66",
  3451 => x"87c2ec49",
  3452 => x"49c086c8",
  3453 => x"ce87c7eb",
  3454 => x"cdef87e8",
  3455 => x"02987087",
  3456 => x"c087dfce",
  3457 => x"496697e5",
  3458 => x"e6c031d0",
  3459 => x"c84a6697",
  3460 => x"c0b17232",
  3461 => x"4a6697e7",
  3462 => x"c74d71b1",
  3463 => x"9dffffff",
  3464 => x"6697e8c0",
  3465 => x"87c8c002",
  3466 => x"a6e4c048",
  3467 => x"87c7c058",
  3468 => x"48a6e0c0",
  3469 => x"7578c0c4",
  3470 => x"87ffe549",
  3471 => x"58eff1c4",
  3472 => x"48daf1c4",
  3473 => x"f1c478c0",
  3474 => x"f1c45df3",
  3475 => x"e0c048f3",
  3476 => x"49757866",
  3477 => x"bfeacbc4",
  3478 => x"f6cbc489",
  3479 => x"cbc491bf",
  3480 => x"7181bfe6",
  3481 => x"fecbc41e",
  3482 => x"c3d4fd49",
  3483 => x"c486c487",
  3484 => x"c048fff1",
  3485 => x"e9f1c478",
  3486 => x"c450c148",
  3487 => x"c248def1",
  3488 => x"87decc50",
  3489 => x"6697e8c0",
  3490 => x"87c9c002",
  3491 => x"48e8f1c4",
  3492 => x"cdcc50c1",
  3493 => x"e849c087",
  3494 => x"c5cc87e4",
  3495 => x"87eaec87",
  3496 => x"cb029870",
  3497 => x"edc087fc",
  3498 => x"48496697",
  3499 => x"c098c0c3",
  3500 => x"7058a6e4",
  3501 => x"dcc00298",
  3502 => x"c0c14887",
  3503 => x"a6e4c088",
  3504 => x"02987058",
  3505 => x"4887e9c0",
  3506 => x"c088c0c1",
  3507 => x"7058a6e4",
  3508 => x"c7c10298",
  3509 => x"97e7c087",
  3510 => x"31d04966",
  3511 => x"6697e8c0",
  3512 => x"7232c84a",
  3513 => x"97e9c0b1",
  3514 => x"714d4a66",
  3515 => x"87f9c0b5",
  3516 => x"6697e8c0",
  3517 => x"87f4e549",
  3518 => x"c01e4970",
  3519 => x"496697eb",
  3520 => x"7087e9e5",
  3521 => x"eec01e49",
  3522 => x"e5496697",
  3523 => x"4a7087de",
  3524 => x"cbc5ff49",
  3525 => x"7086c887",
  3526 => x"87cdc04d",
  3527 => x"6697e6c0",
  3528 => x"87e0e549",
  3529 => x"bfeacbc4",
  3530 => x"daf1c44d",
  3531 => x"c478c048",
  3532 => x"755df3f1",
  3533 => x"87c3e249",
  3534 => x"58eff1c4",
  3535 => x"5dc7f2c4",
  3536 => x"48c7f2c4",
  3537 => x"bfdacbc4",
  3538 => x"cff2c478",
  3539 => x"97e5c048",
  3540 => x"f2c45066",
  3541 => x"78c148cb",
  3542 => x"97cff2c4",
  3543 => x"059949bf",
  3544 => x"c487c9c0",
  3545 => x"c448def1",
  3546 => x"87c6c050",
  3547 => x"48def1c4",
  3548 => x"49c050c3",
  3549 => x"c887ede5",
  3550 => x"cde987e8",
  3551 => x"02987087",
  3552 => x"c087dfc8",
  3553 => x"496697ed",
  3554 => x"98c0c348",
  3555 => x"58a6e4c0",
  3556 => x"c0029870",
  3557 => x"c14887dc",
  3558 => x"e4c088c0",
  3559 => x"987058a6",
  3560 => x"87e9c002",
  3561 => x"88c0c148",
  3562 => x"58a6e4c0",
  3563 => x"c1029870",
  3564 => x"e7c087c7",
  3565 => x"d0496697",
  3566 => x"97e8c031",
  3567 => x"32c84a66",
  3568 => x"e9c0b172",
  3569 => x"4d4a6697",
  3570 => x"eec1b571",
  3571 => x"97e8c087",
  3572 => x"d7e24966",
  3573 => x"1e497087",
  3574 => x"6697ebc0",
  3575 => x"87cce249",
  3576 => x"c01e4970",
  3577 => x"496697ee",
  3578 => x"7087c1e2",
  3579 => x"c1ff494a",
  3580 => x"86c887ee",
  3581 => x"c2c14d70",
  3582 => x"97e6c087",
  3583 => x"ebe14966",
  3584 => x"48497087",
  3585 => x"58a6e4c0",
  3586 => x"c0059870",
  3587 => x"e0c087c6",
  3588 => x"78c148a6",
  3589 => x"4866e0c0",
  3590 => x"bfdecbc4",
  3591 => x"c006a8b7",
  3592 => x"e0c087cc",
  3593 => x"cbc448a6",
  3594 => x"c078bfda",
  3595 => x"e0c087c9",
  3596 => x"cbc448a6",
  3597 => x"c078bfee",
  3598 => x"c44d66e0",
  3599 => x"c048cff2",
  3600 => x"506697e5",
  3601 => x"5dcbf2c4",
  3602 => x"97cff2c4",
  3603 => x"059949bf",
  3604 => x"c487c9c0",
  3605 => x"c048def1",
  3606 => x"87c6c050",
  3607 => x"48def1c4",
  3608 => x"f2c450c3",
  3609 => x"49bf97cf",
  3610 => x"c402a9c2",
  3611 => x"49c087f4",
  3612 => x"c487cbe1",
  3613 => x"d1e587ec",
  3614 => x"02987087",
  3615 => x"c487e3c4",
  3616 => x"c448def1",
  3617 => x"e049c050",
  3618 => x"d5c487f4",
  3619 => x"87fae487",
  3620 => x"c4029870",
  3621 => x"f1c487cc",
  3622 => x"c448bfef",
  3623 => x"88bfeacb",
  3624 => x"58a6e4c0",
  3625 => x"c17e97ca",
  3626 => x"c0c248a6",
  3627 => x"def1c450",
  3628 => x"c048bf97",
  3629 => x"c458a6f7",
  3630 => x"c9c005a8",
  3631 => x"a6f3c087",
  3632 => x"c078c248",
  3633 => x"f3c087e1",
  3634 => x"a8c34866",
  3635 => x"87c9c005",
  3636 => x"48a6f7c0",
  3637 => x"c6c078c0",
  3638 => x"a6f7c087",
  3639 => x"c078c348",
  3640 => x"c048a6f3",
  3641 => x"c27866f7",
  3642 => x"f3c048a6",
  3643 => x"50c05066",
  3644 => x"bfebf1c4",
  3645 => x"ff81c149",
  3646 => x"c487fcdc",
  3647 => x"c45008a6",
  3648 => x"49bfebf1",
  3649 => x"87efdcff",
  3650 => x"5008a6c5",
  3651 => x"4ba6f0c0",
  3652 => x"66e4c01e",
  3653 => x"f7fbfe49",
  3654 => x"97f4c087",
  3655 => x"dcff4966",
  3656 => x"a6ca87d5",
  3657 => x"f5c05008",
  3658 => x"ff496697",
  3659 => x"cb87c8dc",
  3660 => x"c05008a6",
  3661 => x"496697f6",
  3662 => x"87fbdbff",
  3663 => x"5008a6cc",
  3664 => x"f1c41e73",
  3665 => x"fe49bfef",
  3666 => x"c087c5fb",
  3667 => x"496697f8",
  3668 => x"87e3dbff",
  3669 => x"5008a6d1",
  3670 => x"6697f9c0",
  3671 => x"d6dbff49",
  3672 => x"08a6d287",
  3673 => x"97fac050",
  3674 => x"dbff4966",
  3675 => x"a6d387c9",
  3676 => x"1ec15008",
  3677 => x"a6d21eca",
  3678 => x"f5ddff49",
  3679 => x"c086d087",
  3680 => x"f9dcff49",
  3681 => x"87dac087",
  3682 => x"c01e1ec0",
  3683 => x"49c51ee0",
  3684 => x"87d5dcff",
  3685 => x"f1c486cc",
  3686 => x"78c048e4",
  3687 => x"dcff49c1",
  3688 => x"c4ff87dc",
  3689 => x"fbdaff8e",
  3690 => x"86f41e87",
  3691 => x"c848d0ff",
  3692 => x"d4ff78c5",
  3693 => x"78e3c148",
  3694 => x"d4ff4ac0",
  3695 => x"7678c048",
  3696 => x"68817249",
  3697 => x"ca82c151",
  3698 => x"ed04aab7",
  3699 => x"48d0ff87",
  3700 => x"8ef478c4",
  3701 => x"c41e4f26",
  3702 => x"c148e9f1",
  3703 => x"1e4f2650",
  3704 => x"48daf1c4",
  3705 => x"f1c478c0",
  3706 => x"40c048eb",
  3707 => x"f7f1c478",
  3708 => x"c478c048",
  3709 => x"c148dff1",
  3710 => x"c6ccc450",
  3711 => x"87c402bf",
  3712 => x"87c249c0",
  3713 => x"f1c449c1",
  3714 => x"c45997e2",
  3715 => x"c048fbf1",
  3716 => x"f1c47840",
  3717 => x"40c048e4",
  3718 => x"f2c45050",
  3719 => x"40c048c3",
  3720 => x"cff2c478",
  3721 => x"9f50c048",
  3722 => x"eaf1c478",
  3723 => x"2650c148",
  3724 => x"1e731e4f",
  3725 => x"c848d0ff",
  3726 => x"d4ff78c5",
  3727 => x"78e0c148",
  3728 => x"ffc34968",
  3729 => x"48d0ff99",
  3730 => x"4b7178c4",
  3731 => x"0299c149",
  3732 => x"dfe687c3",
  3733 => x"c2497387",
  3734 => x"87c30299",
  3735 => x"7387cafd",
  3736 => x"0299c449",
  3737 => x"edfd87c3",
  3738 => x"c8497387",
  3739 => x"87d60299",
  3740 => x"ff87ecfd",
  3741 => x"c5c848d0",
  3742 => x"48d4ff78",
  3743 => x"c078e6c1",
  3744 => x"48d0ff78",
  3745 => x"497378c4",
  3746 => x"f1c499d0",
  3747 => x"ff5997ee",
  3748 => x"c487dedd",
  3749 => x"02bfe4f1",
  3750 => x"f1c487d7",
  3751 => x"d005bfda",
  3752 => x"d0f2c487",
  3753 => x"ff49bf9f",
  3754 => x"c487d3d8",
  3755 => x"c048e4f1",
  3756 => x"e8f1c478",
  3757 => x"d902bf97",
  3758 => x"48d0ff87",
  3759 => x"ff78c5c8",
  3760 => x"e5c148d4",
  3761 => x"ff78c078",
  3762 => x"78c448d0",
  3763 => x"48e8f1c4",
  3764 => x"d6ff50c0",
  3765 => x"000087d2",
  3766 => x"711e0000",
  3767 => x"bfc8ff4a",
  3768 => x"48a17249",
  3769 => x"ff1e4f26",
  3770 => x"fe89bfc8",
  3771 => x"c0c0c0c0",
  3772 => x"c401a9c0",
  3773 => x"c24ac087",
  3774 => x"724ac187",
  3775 => x"0e4f2648",
  3776 => x"5d5c5b5e",
  3777 => x"ff4b710e",
  3778 => x"66d04cd4",
  3779 => x"d678c048",
  3780 => x"dfcffe49",
  3781 => x"7cffc387",
  3782 => x"ffc3496c",
  3783 => x"494d7199",
  3784 => x"c199f0c3",
  3785 => x"cb05a9e0",
  3786 => x"7cffc387",
  3787 => x"98c3486c",
  3788 => x"780866d0",
  3789 => x"6c7cffc3",
  3790 => x"31c8494a",
  3791 => x"6c7cffc3",
  3792 => x"72b2714a",
  3793 => x"c331c849",
  3794 => x"4a6c7cff",
  3795 => x"4972b271",
  3796 => x"ffc331c8",
  3797 => x"714a6c7c",
  3798 => x"48d0ffb2",
  3799 => x"7378e0c0",
  3800 => x"87c2029b",
  3801 => x"48757b72",
  3802 => x"4c264d26",
  3803 => x"4f264b26",
  3804 => x"0e4f261e",
  3805 => x"0e5c5b5e",
  3806 => x"1e7686f8",
  3807 => x"fd49a6c8",
  3808 => x"86c487fd",
  3809 => x"486e4b70",
  3810 => x"c201a8c0",
  3811 => x"4a7387f0",
  3812 => x"c19af0c3",
  3813 => x"c702aad0",
  3814 => x"aae0c187",
  3815 => x"87dec205",
  3816 => x"99c84973",
  3817 => x"ff87c302",
  3818 => x"4c7387c6",
  3819 => x"acc29cc3",
  3820 => x"87c2c105",
  3821 => x"c94966c4",
  3822 => x"c41e7131",
  3823 => x"92d44a66",
  3824 => x"49d2f2c4",
  3825 => x"fefc8172",
  3826 => x"49d887e6",
  3827 => x"87e4ccfe",
  3828 => x"c31ec0c8",
  3829 => x"fc49cafa",
  3830 => x"ff87ffda",
  3831 => x"e0c048d0",
  3832 => x"cafac378",
  3833 => x"4a66cc1e",
  3834 => x"f2c492d4",
  3835 => x"817249d2",
  3836 => x"87f9fcfc",
  3837 => x"acc186cc",
  3838 => x"87c2c105",
  3839 => x"c94966c4",
  3840 => x"c41e7131",
  3841 => x"92d44a66",
  3842 => x"49d2f2c4",
  3843 => x"fdfc8172",
  3844 => x"fac387de",
  3845 => x"66c81eca",
  3846 => x"c492d44a",
  3847 => x"7249d2f2",
  3848 => x"c5fbfc81",
  3849 => x"fe49d787",
  3850 => x"c887c9cb",
  3851 => x"fac31ec0",
  3852 => x"d9fc49ca",
  3853 => x"86cc87ce",
  3854 => x"c048d0ff",
  3855 => x"8ef878e0",
  3856 => x"0e87e7fc",
  3857 => x"5d5c5b5e",
  3858 => x"4d711e0e",
  3859 => x"d44cd4ff",
  3860 => x"c3487e66",
  3861 => x"c506a8b7",
  3862 => x"c148c087",
  3863 => x"497587e2",
  3864 => x"87cad1fd",
  3865 => x"66c41e75",
  3866 => x"c493d44b",
  3867 => x"7383d2f2",
  3868 => x"d9f6fc49",
  3869 => x"6b83c887",
  3870 => x"48d0ff4b",
  3871 => x"dd78e1c8",
  3872 => x"c349737c",
  3873 => x"7c7199ff",
  3874 => x"b7c84973",
  3875 => x"99ffc329",
  3876 => x"49737c71",
  3877 => x"c329b7d0",
  3878 => x"7c7199ff",
  3879 => x"b7d84973",
  3880 => x"c07c7129",
  3881 => x"7c7c7c7c",
  3882 => x"7c7c7c7c",
  3883 => x"7c7c7c7c",
  3884 => x"c478e0c0",
  3885 => x"49dc1e66",
  3886 => x"87ddc9fe",
  3887 => x"487386c8",
  3888 => x"87e4fa26",
  3889 => x"5c5b5e0e",
  3890 => x"711e0e5d",
  3891 => x"4bd4ff7e",
  3892 => x"f2c41e6e",
  3893 => x"f4fc49e6",
  3894 => x"86c487f4",
  3895 => x"029d4d70",
  3896 => x"c487c3c3",
  3897 => x"4cbfeef2",
  3898 => x"cffd496e",
  3899 => x"d0ff87c0",
  3900 => x"78c5c848",
  3901 => x"c07bd6c1",
  3902 => x"c17b154a",
  3903 => x"b7e0c082",
  3904 => x"87f504aa",
  3905 => x"c448d0ff",
  3906 => x"78c5c878",
  3907 => x"c17bd3c1",
  3908 => x"7478c47b",
  3909 => x"fcc1029c",
  3910 => x"cafac387",
  3911 => x"4dc0c87e",
  3912 => x"acb7c08c",
  3913 => x"c887c603",
  3914 => x"c04da4c0",
  3915 => x"fbc6c44c",
  3916 => x"d049bf97",
  3917 => x"87d20299",
  3918 => x"f2c41ec0",
  3919 => x"f6fc49e6",
  3920 => x"86c487e8",
  3921 => x"c04a4970",
  3922 => x"fac387ef",
  3923 => x"f2c41eca",
  3924 => x"f6fc49e6",
  3925 => x"86c487d4",
  3926 => x"ff4a4970",
  3927 => x"c5c848d0",
  3928 => x"7bd4c178",
  3929 => x"7bbf976e",
  3930 => x"80c1486e",
  3931 => x"8dc17e70",
  3932 => x"87f0ff05",
  3933 => x"c448d0ff",
  3934 => x"059a7278",
  3935 => x"48c087c5",
  3936 => x"c187e5c0",
  3937 => x"e6f2c41e",
  3938 => x"fcf3fc49",
  3939 => x"7486c487",
  3940 => x"c4fe059c",
  3941 => x"48d0ff87",
  3942 => x"c178c5c8",
  3943 => x"7bc07bd3",
  3944 => x"48c178c4",
  3945 => x"48c087c2",
  3946 => x"264d2626",
  3947 => x"264b264c",
  3948 => x"5b5e0e4f",
  3949 => x"4b710e5c",
  3950 => x"dd0266cc",
  3951 => x"f0c04c87",
  3952 => x"87dd028c",
  3953 => x"8ac14a74",
  3954 => x"8a87d602",
  3955 => x"8a87d202",
  3956 => x"d087ce02",
  3957 => x"87db028a",
  3958 => x"497387df",
  3959 => x"d887e5fb",
  3960 => x"c01e7487",
  3961 => x"87dbf949",
  3962 => x"49731e74",
  3963 => x"c887d4f9",
  3964 => x"7387c686",
  3965 => x"ccd0fd49",
  3966 => x"87effe87",
  3967 => x"f9c31e00",
  3968 => x"c149bfcb",
  3969 => x"cff9c3b9",
  3970 => x"48d4ff59",
  3971 => x"ff78ffc3",
  3972 => x"e1c848d0",
  3973 => x"48d4ff78",
  3974 => x"31c478c1",
  3975 => x"d0ff7871",
  3976 => x"78e0c048",
  3977 => x"c31e4f26",
  3978 => x"c41efff8",
  3979 => x"fc49e6f2",
  3980 => x"c487dbef",
  3981 => x"02987086",
  3982 => x"c0ff87c3",
  3983 => x"314f2687",
  3984 => x"5a484b35",
  3985 => x"43202020",
  3986 => x"00004746",
  3987 => x"1a000000",
  3988 => x"1112589f",
  3989 => x"1c1b1d14",
  3990 => x"5aa74a23",
  3991 => x"f5949159",
  3992 => x"f5f4ebf2",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
